magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_s >>
rect 8516 8522 9286 10772
<< dnwell >>
rect 8516 8522 9286 10772
<< nwell >>
rect 8422 10452 9358 10738
rect 8422 8772 8708 10452
rect 9072 8772 9358 10452
rect 8422 8486 9358 8772
<< pwell >>
rect 9473 7000 9486 7008
rect 9473 6908 9486 6910
rect 10082 6740 10118 6868
rect 10184 6738 10234 6882
rect 10886 6800 10906 6902
rect 4158 4578 4288 4712
<< nsubdiff >>
rect 8459 10681 9321 10701
rect 8459 10647 8539 10681
rect 9241 10647 9321 10681
rect 8459 10627 9321 10647
rect 8459 10621 8533 10627
rect 8459 8603 8479 10621
rect 8513 8603 8533 10621
rect 8459 8597 8533 8603
rect 9247 10621 9321 10627
rect 9247 8603 9267 10621
rect 9301 8603 9321 10621
rect 9247 8597 9321 8603
rect 8459 8577 9321 8597
rect 8459 8543 8539 8577
rect 9241 8543 9321 8577
rect 8459 8523 9321 8543
<< nsubdiffcont >>
rect 8539 10647 9241 10681
rect 8479 8603 8513 10621
rect 9267 8603 9301 10621
rect 8539 8543 9241 8577
<< locali >>
rect 8479 10647 8539 10681
rect 9241 10647 9301 10681
rect 8479 10621 8513 10647
rect 6568 10108 6718 10170
rect 4138 9548 4732 9696
rect 4142 5642 4298 9548
rect 6590 9056 6736 9130
rect 9267 10621 9301 10647
rect 8479 8577 8513 8603
rect 11982 8758 14642 8900
rect 9267 8577 9301 8603
rect 8479 8543 8539 8577
rect 9241 8543 9301 8577
rect 8114 8362 8514 8384
rect 8672 8362 8698 8384
rect 8114 8260 8698 8362
rect 6614 7942 6760 8016
rect 14326 7808 14420 7884
rect 8062 6968 8222 7142
rect 8500 6532 8634 6850
rect 14540 6766 14636 8758
rect 11506 6714 14642 6766
rect 11344 6678 14642 6714
rect 7792 6144 7944 6218
rect 4596 5642 4710 6002
rect 4142 5534 4710 5642
rect 8706 5774 9052 5884
rect 4148 5526 4710 5534
rect 4596 4676 4710 5526
rect 4596 4570 5878 4676
rect 4596 4538 4710 4570
rect 4458 4502 4710 4538
<< viali >>
rect 8098 8866 8148 8958
rect 9182 8910 9228 9096
rect 10356 9560 10406 9706
rect 9260 8930 9267 9078
rect 9267 8930 9301 9078
rect 9301 8930 9322 9078
rect 8890 8577 8988 8582
rect 8890 8543 8988 8577
rect 8890 8536 8988 8543
rect 7878 8178 7948 8286
rect 11280 7108 11336 7150
rect 10918 7050 10954 7088
rect 10122 6978 10156 7012
rect 11084 6976 11146 7024
rect 10010 6904 10066 6944
rect 10344 6480 10484 6518
rect 5442 5626 5552 5838
rect 9028 5660 9206 5724
rect 4288 4738 4330 4776
rect 4430 4740 4486 4780
<< metal1 >>
rect 6772 10722 6782 10936
rect 6998 10722 7008 10936
rect 7602 10682 8112 10698
rect 7602 10590 9132 10682
rect 7602 10570 8112 10590
rect 5544 10482 6562 10496
rect 5484 10408 6562 10482
rect 5484 10378 5550 10408
rect 4830 9932 4840 10346
rect 5098 9932 5108 10346
rect 5484 9980 5494 10378
rect 5556 9980 5566 10378
rect 6550 9984 6560 10378
rect 6614 9984 6624 10378
rect 6662 10120 6672 10262
rect 6732 10120 6742 10262
rect 5484 9950 5550 9980
rect 5484 9862 6602 9950
rect 7576 9868 7586 10024
rect 7638 9868 7648 10024
rect 7778 9866 7788 10022
rect 7840 9866 7850 10022
rect 7966 9872 7976 10028
rect 8028 9872 8038 10028
rect 4826 9682 4836 9708
rect 4794 9294 4836 9682
rect 5094 9294 5104 9708
rect 5886 9692 6136 9862
rect 6832 9692 6930 9698
rect 5886 9592 6938 9692
rect 5510 9392 5592 9398
rect 5508 9316 6576 9392
rect 4346 8764 4574 8780
rect 4794 8764 5088 9294
rect 5510 9244 5592 9316
rect 5506 9002 5516 9244
rect 5570 9002 5592 9244
rect 6832 9180 6930 9592
rect 5510 8856 5592 9002
rect 6558 8998 6568 9180
rect 6646 9172 6978 9180
rect 6646 9024 6700 9172
rect 6758 9024 6978 9172
rect 6646 8998 6978 9024
rect 6574 8996 6978 8998
rect 6832 8992 6930 8996
rect 5950 8856 6146 8874
rect 5510 8792 6578 8856
rect 7676 8834 7686 8990
rect 7738 8834 7748 8990
rect 7874 8828 7884 8984
rect 7936 8828 7946 8984
rect 8092 8966 8154 8970
rect 8088 8872 8098 8966
rect 8154 8872 8164 8966
rect 8092 8866 8098 8872
rect 8148 8866 8154 8872
rect 8092 8854 8154 8866
rect 5510 8766 5592 8792
rect 4346 8552 5088 8764
rect 5950 8730 6146 8792
rect 5954 8604 6144 8730
rect 7494 8706 8004 8708
rect 8256 8706 8336 10590
rect 8648 9868 8658 10078
rect 8734 9868 8744 10078
rect 8846 9864 8856 10074
rect 8932 9864 8942 10074
rect 9036 9862 9046 10072
rect 9122 10032 9132 10072
rect 9122 9864 9514 10032
rect 9122 9862 9132 9864
rect 9400 9814 9514 9864
rect 9400 9812 9864 9814
rect 9400 9740 10284 9812
rect 9400 9738 9864 9740
rect 9400 9716 9536 9738
rect 9434 9276 9536 9716
rect 10350 9706 10412 9718
rect 9728 9568 9738 9672
rect 9812 9568 9822 9672
rect 9936 9562 9946 9666
rect 10000 9562 10010 9666
rect 10122 9560 10132 9664
rect 10186 9560 10196 9664
rect 10350 9660 10356 9706
rect 10406 9660 10412 9706
rect 10346 9560 10356 9660
rect 10424 9560 10434 9660
rect 10350 9548 10412 9560
rect 11616 9444 11626 9866
rect 11874 9444 11884 9866
rect 9838 9332 9848 9436
rect 9902 9332 9912 9436
rect 10028 9330 10038 9434
rect 10092 9330 10102 9434
rect 10220 9334 10230 9438
rect 10284 9334 10294 9438
rect 9434 9274 9986 9276
rect 9434 9202 10276 9274
rect 9434 9200 9986 9202
rect 9490 9186 9986 9200
rect 9176 9096 9234 9108
rect 9176 9088 9182 9096
rect 9228 9090 9300 9096
rect 9228 9088 9328 9090
rect 8550 8968 8620 8980
rect 8756 8916 8766 9072
rect 8818 8916 8828 9072
rect 8948 8922 8958 9078
rect 9010 8922 9020 9078
rect 9158 8922 9168 9088
rect 9240 9078 9328 9088
rect 9240 8930 9260 9078
rect 9322 8930 9332 9078
rect 9240 8922 9328 8930
rect 8962 8888 8970 8922
rect 9176 8910 9182 8922
rect 9228 8918 9328 8922
rect 9228 8914 9300 8918
rect 9228 8910 9234 8914
rect 9176 8898 9234 8910
rect 8964 8876 8970 8888
rect 11596 8812 11606 9218
rect 11888 8812 11898 9218
rect 8550 8796 8620 8808
rect 9068 8792 9072 8810
rect 8646 8706 9156 8718
rect 7494 8622 9156 8706
rect 7494 8620 9036 8622
rect 6862 8604 6972 8606
rect 4346 7732 4574 8552
rect 4794 8550 5088 8552
rect 5946 8518 6972 8604
rect 7494 8580 8004 8620
rect 8646 8590 9036 8620
rect 8878 8582 9000 8588
rect 6062 8516 6972 8518
rect 5542 8274 5606 8276
rect 5542 8206 6600 8274
rect 5542 8174 5606 8206
rect 5528 7776 5538 8174
rect 5600 7776 5610 8174
rect 6588 8116 6698 8178
rect 6588 7900 6600 8116
rect 6664 8100 6698 8116
rect 6664 8052 6694 8100
rect 6862 8052 6972 8516
rect 6664 7924 6726 8052
rect 6786 7924 6972 8052
rect 6664 7922 6972 7924
rect 6664 7900 6694 7922
rect 6584 7782 6690 7900
rect 5542 7736 5606 7776
rect 4346 7528 4364 7732
rect 4354 7526 4364 7528
rect 4558 7726 4574 7732
rect 5160 7732 5654 7736
rect 5160 7728 6592 7732
rect 4558 7526 4900 7726
rect 4636 7158 4900 7526
rect 5154 7678 6592 7728
rect 5154 7662 5654 7678
rect 7564 7676 7818 8580
rect 8878 8536 8890 8582
rect 8988 8536 9000 8582
rect 9024 8566 9036 8590
rect 9130 8590 9156 8622
rect 9130 8566 9142 8590
rect 9024 8560 9142 8566
rect 8878 8530 9000 8536
rect 7872 8286 7954 8298
rect 7994 8288 8056 8338
rect 7868 8178 7878 8286
rect 7948 8178 7958 8286
rect 7994 8210 8068 8288
rect 8728 8210 8778 8296
rect 7994 8208 8802 8210
rect 8924 8208 8980 8530
rect 7996 8200 9022 8208
rect 7872 8166 7954 8178
rect 7996 8160 8348 8200
rect 8008 8154 8348 8160
rect 8338 8146 8348 8154
rect 8484 8162 9022 8200
rect 8484 8154 8802 8162
rect 8924 8158 8980 8162
rect 8484 8146 8494 8154
rect 9206 7762 9216 7972
rect 9278 7762 9288 7972
rect 14276 7778 14286 7964
rect 14338 7778 14348 7964
rect 7558 7670 8570 7676
rect 4616 6724 4626 7158
rect 4902 6724 4912 7158
rect 4636 6722 4900 6724
rect 4078 6402 4544 6404
rect 4616 6402 4626 6488
rect 3574 6398 3848 6400
rect 4078 6398 4626 6402
rect 3574 6116 4626 6398
rect 3574 6110 4110 6116
rect 4458 6110 4626 6116
rect 3574 4788 3848 6110
rect 4616 6054 4626 6110
rect 4902 6402 4912 6488
rect 4902 6110 4924 6402
rect 4902 6054 4912 6110
rect 5154 5842 5334 7662
rect 7548 7570 8570 7670
rect 7548 7530 7802 7570
rect 7548 7408 7818 7530
rect 8462 7492 8564 7570
rect 7564 7282 7818 7408
rect 6500 7194 6968 7228
rect 5732 7112 6968 7194
rect 5582 6624 5592 7080
rect 5650 6624 5660 7080
rect 5774 6620 5784 7076
rect 5842 6620 5852 7076
rect 5968 6626 5978 7082
rect 6036 6626 6046 7082
rect 6160 6624 6170 7080
rect 6228 6624 6238 7080
rect 6354 6624 6364 7080
rect 6422 6624 6432 7080
rect 6546 6620 6556 7076
rect 6614 6620 6624 7076
rect 5436 5842 5558 5850
rect 5160 5834 5362 5842
rect 5436 5838 5466 5842
rect 5532 5838 5558 5842
rect 5436 5834 5442 5838
rect 5160 5650 5442 5834
rect 5160 5646 5362 5650
rect 5436 5626 5442 5650
rect 5552 5626 5558 5838
rect 5678 5842 5688 5966
rect 5746 5842 5756 5966
rect 5678 5834 5756 5842
rect 5436 5614 5558 5626
rect 5678 5510 5688 5650
rect 5746 5510 5756 5650
rect 5872 5520 5882 5976
rect 5940 5520 5950 5976
rect 6064 5518 6074 5974
rect 6132 5518 6142 5974
rect 6256 5504 6266 5960
rect 6324 5504 6334 5960
rect 6448 5504 6458 5960
rect 6516 5504 6526 5960
rect 6886 5454 6968 7112
rect 7564 7074 7574 7282
rect 7756 7160 7818 7282
rect 7916 7280 7926 7438
rect 8020 7280 8030 7438
rect 8462 7424 9092 7492
rect 8468 7420 9092 7424
rect 8398 7272 8408 7378
rect 8464 7272 8474 7378
rect 8590 7270 8600 7376
rect 8656 7270 8666 7376
rect 8792 7268 8802 7374
rect 8858 7268 8868 7374
rect 7756 7074 7816 7160
rect 7564 6914 7816 7074
rect 8048 6976 8058 7134
rect 8152 6976 8162 7134
rect 8504 7034 8514 7140
rect 8570 7034 8580 7140
rect 8692 7036 8702 7142
rect 8758 7036 8768 7142
rect 8882 7024 8892 7148
rect 8956 7024 8966 7148
rect 9002 6962 9092 7420
rect 9236 7346 9528 7724
rect 9234 7244 9266 7346
rect 9412 7244 9528 7346
rect 9234 7200 9528 7244
rect 9236 7190 9528 7200
rect 9240 7180 9436 7190
rect 9950 7186 9960 7276
rect 10044 7186 10054 7276
rect 10862 7242 10872 7326
rect 10970 7242 10980 7326
rect 7558 6910 7956 6914
rect 7558 6906 8238 6910
rect 8372 6906 9092 6962
rect 9244 6978 9436 7180
rect 11630 7156 11830 7290
rect 11268 7150 11832 7156
rect 11268 7108 11280 7150
rect 11336 7108 11832 7150
rect 11268 7102 11348 7108
rect 10912 7098 10960 7100
rect 10900 7030 10910 7098
rect 10970 7030 10980 7098
rect 11630 7092 11830 7108
rect 11072 7024 11158 7030
rect 10122 7018 10350 7022
rect 10110 7012 10350 7018
rect 10110 6978 10122 7012
rect 10156 6996 10350 7012
rect 11072 6996 11084 7024
rect 10156 6984 11084 6996
rect 10156 6978 10228 6984
rect 9244 6958 9494 6978
rect 10110 6972 10228 6978
rect 10296 6976 11084 6984
rect 11146 6976 11158 7024
rect 10296 6970 11158 6976
rect 10296 6968 11150 6970
rect 9244 6950 9896 6958
rect 9244 6944 10078 6950
rect 9244 6912 10010 6944
rect 7558 6902 9092 6906
rect 9216 6904 10010 6912
rect 10066 6904 10078 6944
rect 7558 6898 9088 6902
rect 7558 6850 8438 6898
rect 8766 6896 8980 6898
rect 9216 6896 10078 6904
rect 7558 6840 8404 6850
rect 9216 6842 9896 6896
rect 7558 6838 8238 6840
rect 7840 6834 8238 6838
rect 7960 6714 7970 6792
rect 8114 6714 8124 6792
rect 9216 6748 9522 6842
rect 10856 6772 10866 6790
rect 9012 6662 9552 6748
rect 9010 6580 9552 6662
rect 9938 6724 10070 6760
rect 10824 6724 10866 6772
rect 9938 6660 9952 6724
rect 10044 6660 10070 6724
rect 10856 6686 10866 6724
rect 10996 6686 11006 6790
rect 9952 6640 9962 6660
rect 7344 6502 8634 6504
rect 9010 6502 9092 6580
rect 9428 6566 9500 6580
rect 10334 6524 10344 6548
rect 7344 6420 9092 6502
rect 10332 6480 10344 6524
rect 10482 6524 10492 6548
rect 10482 6518 10496 6524
rect 10484 6480 10496 6518
rect 10332 6474 10496 6480
rect 10434 6434 12558 6444
rect 7344 6418 9034 6420
rect 7344 6416 8634 6418
rect 7346 6350 7454 6416
rect 7346 6302 7782 6350
rect 7348 6284 7782 6302
rect 7348 6026 7452 6284
rect 8278 6256 8288 6382
rect 8342 6256 8352 6382
rect 8470 6256 8480 6382
rect 8534 6256 8544 6382
rect 9634 6362 12558 6434
rect 9634 6358 9714 6362
rect 8674 6282 8684 6354
rect 8760 6282 8770 6354
rect 9586 6332 9714 6358
rect 7784 6166 7794 6234
rect 7860 6166 7870 6234
rect 9586 6176 9698 6332
rect 9580 6174 9728 6176
rect 8958 6170 9728 6174
rect 7502 6134 7588 6142
rect 7502 6058 7512 6134
rect 7578 6058 7588 6134
rect 8168 6134 8254 6142
rect 8168 6058 8178 6134
rect 8244 6058 8254 6134
rect 8366 6132 8452 6140
rect 8366 6056 8376 6132
rect 8442 6056 8452 6132
rect 8562 6138 8648 6142
rect 8948 6138 9728 6170
rect 8562 6134 9728 6138
rect 8562 6058 8572 6134
rect 8638 6098 9728 6134
rect 8638 6094 9414 6098
rect 8638 6058 9042 6094
rect 8578 6046 9042 6058
rect 8948 6028 9040 6046
rect 7348 6002 7458 6026
rect 7348 5946 7798 6002
rect 7350 5944 7798 5946
rect 7350 5758 7458 5944
rect 8960 5838 9024 6028
rect 9368 6000 9378 6062
rect 9444 6000 9454 6062
rect 9580 5960 9728 6098
rect 9104 5868 9114 5932
rect 9166 5868 9176 5932
rect 9582 5892 9728 5960
rect 8944 5758 9400 5838
rect 7350 5664 8738 5758
rect 9016 5726 9218 5730
rect 7350 5654 7458 5664
rect 9014 5662 9024 5726
rect 9202 5724 9218 5726
rect 9016 5660 9028 5662
rect 9206 5660 9218 5724
rect 9016 5654 9218 5660
rect 5626 5448 6276 5454
rect 6358 5448 6968 5454
rect 5626 5380 6968 5448
rect 6254 5192 6336 5380
rect 6366 5370 6968 5380
rect 7874 5192 7904 5398
rect 8122 5192 8132 5398
rect 4222 5100 4232 5124
rect 4014 5024 4232 5100
rect 4306 5100 4316 5124
rect 4306 5024 4360 5100
rect 4014 5016 4360 5024
rect 4598 5088 6338 5192
rect 4598 4790 4678 5088
rect 6254 4968 6336 5088
rect 5964 4916 6336 4968
rect 5964 4900 6356 4916
rect 6024 4804 6034 4860
rect 6092 4804 6102 4860
rect 6136 4806 6146 4862
rect 6204 4806 6214 4862
rect 3566 4776 4354 4788
rect 4430 4786 4680 4790
rect 3566 4738 4288 4776
rect 4330 4738 4354 4776
rect 3566 4712 4354 4738
rect 4418 4780 4680 4786
rect 4418 4740 4430 4780
rect 4486 4774 4680 4780
rect 4486 4740 4682 4774
rect 4418 4734 4682 4740
rect 4434 4730 4682 4734
rect 5916 4684 5926 4740
rect 5984 4684 5994 4740
rect 6274 4642 6356 4900
rect 9580 4700 9728 5892
rect 10062 5882 10072 6126
rect 10162 5882 10172 6126
rect 10398 5876 10408 6120
rect 10584 5888 10594 6140
rect 10678 5888 10688 6140
rect 10914 5876 10924 6120
rect 11100 5872 11110 6124
rect 11194 5872 11204 6124
rect 11428 5890 11438 6134
rect 11618 5864 11628 6116
rect 11712 5864 11722 6116
rect 11944 5868 11954 6112
rect 12130 5864 12140 6116
rect 12224 5864 12234 6116
rect 12642 5878 12652 6130
rect 12736 5878 12746 6130
rect 10332 5122 10408 5188
rect 10330 4924 10340 5122
rect 10416 4924 10426 5122
rect 10836 4932 10846 5142
rect 10950 4932 10960 5142
rect 11360 4918 11370 5128
rect 11474 4918 11484 5128
rect 11864 4928 11874 5138
rect 11978 4928 11988 5138
rect 12382 4932 12392 5142
rect 12496 4932 12506 5142
rect 5944 4560 6356 4642
rect 9544 4616 12570 4700
rect 4070 4552 4314 4556
rect 4070 4476 4230 4552
rect 4220 4474 4230 4476
rect 4304 4474 4314 4552
<< via1 >>
rect 6782 10722 6998 10936
rect 4840 9932 5098 10346
rect 5494 9980 5556 10378
rect 6560 9984 6614 10378
rect 6672 10120 6732 10262
rect 7586 9868 7638 10024
rect 7788 9866 7840 10022
rect 7976 9872 8028 10028
rect 4836 9294 5094 9708
rect 5516 9002 5570 9244
rect 6568 8998 6646 9180
rect 6700 9024 6758 9172
rect 7686 8834 7738 8990
rect 7884 8828 7936 8984
rect 8098 8958 8154 8966
rect 8098 8872 8148 8958
rect 8148 8872 8154 8958
rect 8658 9868 8734 10078
rect 8856 9864 8932 10074
rect 9046 9862 9122 10072
rect 9738 9568 9812 9672
rect 9946 9562 10000 9666
rect 10132 9560 10186 9664
rect 10356 9560 10406 9660
rect 10406 9560 10424 9660
rect 11626 9444 11874 9866
rect 9848 9332 9902 9436
rect 10038 9330 10092 9434
rect 10230 9334 10284 9438
rect 8766 8916 8818 9072
rect 8958 8922 9010 9078
rect 9168 8922 9182 9088
rect 9182 8922 9228 9088
rect 9228 8922 9240 9088
rect 9260 8930 9322 9078
rect 11606 8812 11888 9218
rect 5538 7776 5600 8174
rect 6600 7900 6664 8116
rect 6726 7924 6786 8052
rect 4364 7526 4558 7732
rect 7878 8178 7948 8286
rect 8348 8146 8484 8200
rect 9216 7762 9278 7972
rect 14286 7778 14338 7964
rect 4626 6724 4902 7158
rect 4626 6054 4902 6488
rect 5592 6624 5650 7080
rect 5784 6620 5842 7076
rect 5978 6626 6036 7082
rect 6170 6624 6228 7080
rect 6364 6624 6422 7080
rect 6556 6620 6614 7076
rect 5466 5838 5532 5842
rect 5466 5642 5532 5838
rect 5688 5842 5746 5966
rect 5688 5510 5746 5650
rect 5882 5520 5940 5976
rect 6074 5518 6132 5974
rect 6266 5504 6324 5960
rect 6458 5504 6516 5960
rect 7574 7074 7756 7282
rect 7926 7280 8020 7438
rect 8408 7272 8464 7378
rect 8600 7270 8656 7376
rect 8802 7268 8858 7374
rect 8058 6976 8152 7134
rect 8514 7034 8570 7140
rect 8702 7036 8758 7142
rect 8892 7024 8956 7148
rect 9266 7244 9412 7346
rect 9960 7186 10044 7276
rect 10872 7242 10970 7326
rect 10910 7088 10970 7098
rect 10910 7050 10918 7088
rect 10918 7050 10954 7088
rect 10954 7050 10970 7088
rect 10910 7030 10970 7050
rect 7970 6714 8114 6792
rect 9952 6660 10044 6724
rect 10866 6686 10996 6790
rect 10344 6518 10482 6548
rect 10344 6480 10482 6518
rect 8288 6256 8342 6382
rect 8480 6256 8534 6382
rect 8684 6282 8760 6354
rect 7794 6166 7860 6234
rect 7512 6058 7578 6134
rect 8178 6058 8244 6134
rect 8376 6056 8442 6132
rect 8572 6058 8638 6134
rect 9378 6000 9444 6062
rect 9114 5868 9166 5932
rect 9024 5724 9202 5726
rect 9024 5662 9028 5724
rect 9028 5662 9202 5724
rect 7904 5192 8122 5398
rect 4232 5024 4306 5124
rect 6034 4804 6092 4860
rect 6146 4806 6204 4862
rect 5926 4684 5984 4740
rect 10072 5882 10162 6126
rect 10594 5888 10678 6140
rect 11110 5872 11194 6124
rect 11628 5864 11712 6116
rect 12140 5864 12224 6116
rect 12652 5878 12736 6130
rect 10340 4924 10416 5122
rect 10846 4932 10950 5142
rect 11370 4918 11474 5128
rect 11874 4928 11978 5138
rect 12392 4932 12496 5142
rect 4230 4474 4304 4552
<< metal2 >>
rect 6782 10936 6998 10946
rect 6998 10722 7008 10918
rect 6782 10710 7008 10722
rect 5494 10378 5556 10388
rect 4840 10346 5098 10356
rect 6560 10378 6614 10388
rect 6558 10290 6560 10300
rect 6614 10290 6628 10300
rect 6682 10282 6752 10292
rect 6558 10116 6560 10126
rect 5494 9970 5556 9980
rect 6614 10116 6628 10126
rect 6672 10262 6682 10272
rect 6672 10118 6682 10120
rect 6672 10110 6752 10118
rect 6682 10108 6752 10110
rect 8658 10084 8734 10088
rect 7596 10078 9166 10084
rect 7596 10034 8658 10078
rect 6560 9974 6614 9984
rect 7586 10028 8658 10034
rect 7586 10024 7976 10028
rect 4840 9922 5098 9932
rect 7638 10022 7976 10024
rect 7638 9872 7788 10022
rect 7586 9858 7638 9868
rect 7840 9872 7976 10022
rect 8028 9872 8658 10028
rect 7788 9856 7840 9866
rect 7976 9862 8028 9872
rect 8734 10074 9166 10078
rect 8734 9872 8856 10074
rect 8658 9858 8734 9868
rect 8932 10072 9166 10074
rect 8932 9872 9046 10072
rect 8856 9854 8932 9864
rect 9122 9872 9166 10072
rect 9046 9852 9122 9862
rect 11622 9868 11874 9878
rect 4836 9708 5094 9718
rect 4836 9284 5094 9294
rect 9712 9682 9786 9702
rect 9712 9676 9812 9682
rect 9712 9672 10196 9676
rect 9712 9568 9738 9672
rect 9812 9666 10196 9672
rect 9812 9568 9946 9666
rect 9712 9558 9812 9568
rect 10000 9664 10196 9666
rect 10000 9568 10132 9664
rect 5516 9244 5570 9254
rect 5516 8992 5570 9002
rect 6568 9180 6646 9190
rect 6700 9172 6758 9182
rect 8946 9088 9022 9098
rect 8766 9076 8818 9082
rect 8942 9076 8946 9082
rect 9168 9088 9240 9098
rect 6700 9014 6758 9024
rect 8758 9072 8946 9076
rect 8096 9002 8172 9012
rect 6568 8988 6646 8998
rect 7686 8990 7738 9000
rect 7884 8988 7936 8994
rect 7738 8986 7940 8988
rect 7738 8984 8096 8986
rect 7738 8836 7884 8984
rect 7874 8834 7884 8836
rect 7686 8824 7738 8834
rect 7936 8860 8096 8984
rect 8172 8860 8174 8986
rect 8758 8916 8766 9072
rect 8818 8918 8946 9072
rect 9022 8922 9168 9082
rect 9260 9082 9322 9088
rect 9240 9078 9324 9082
rect 9240 8930 9260 9078
rect 9322 8930 9324 9078
rect 9240 8922 9324 8930
rect 9022 8918 9324 8922
rect 8818 8916 9324 8918
rect 8766 8906 8818 8916
rect 8942 8912 9324 8916
rect 8946 8908 9022 8912
rect 7936 8834 8174 8860
rect 7884 8818 7936 8828
rect 9036 8622 9130 8632
rect 9036 8556 9130 8566
rect 9208 8478 9290 8488
rect 9712 8478 9786 9558
rect 9946 9552 10000 9562
rect 10186 9568 10196 9664
rect 10356 9660 10424 9670
rect 10132 9550 10186 9560
rect 10356 9550 10424 9560
rect 9838 9452 9912 9460
rect 9838 9450 10304 9452
rect 9912 9438 10304 9450
rect 11622 9444 11626 9454
rect 9912 9434 10230 9438
rect 9912 9330 10038 9434
rect 10092 9334 10230 9434
rect 10284 9334 10304 9438
rect 11626 9434 11874 9444
rect 10092 9330 10304 9334
rect 9912 9324 10304 9330
rect 9838 9320 10304 9324
rect 9838 9314 9912 9320
rect 11606 9218 11888 9228
rect 11606 8802 11888 8812
rect 9198 8352 9852 8478
rect 7878 8286 7948 8296
rect 5538 8174 5600 8184
rect 7878 8168 7948 8178
rect 8348 8200 8484 8210
rect 8348 8136 8484 8146
rect 6600 8116 6664 8128
rect 6726 8052 6786 8062
rect 9208 7972 9290 8352
rect 9208 7964 9216 7972
rect 6726 7914 6786 7924
rect 6600 7890 6664 7900
rect 6602 7880 6656 7890
rect 5538 7766 5600 7776
rect 7572 7762 9216 7964
rect 9278 7782 9290 7972
rect 14286 7964 14338 7974
rect 14338 7914 14352 7924
rect 9278 7762 9286 7782
rect 14338 7812 14352 7822
rect 14286 7768 14338 7778
rect 7572 7756 9286 7762
rect 4364 7732 4558 7742
rect 4364 7516 4558 7526
rect 7580 7684 7766 7756
rect 9216 7752 9278 7756
rect 7074 7284 7196 7330
rect 7580 7298 7764 7684
rect 7926 7438 8020 7448
rect 7574 7284 7764 7298
rect 7908 7286 7926 7392
rect 7074 7282 7776 7284
rect 4626 7158 4902 7168
rect 7074 7104 7574 7282
rect 5592 7080 5650 7090
rect 4626 6714 4902 6724
rect 5562 6626 5592 7058
rect 5784 7076 5842 7086
rect 5650 6626 5784 7058
rect 5592 6614 5650 6624
rect 5978 7082 6036 7092
rect 5842 6626 5978 7058
rect 6170 7080 6228 7090
rect 6036 6626 6170 7058
rect 5784 6610 5842 6620
rect 5978 6616 6036 6626
rect 6364 7080 6422 7090
rect 6228 6626 6364 7058
rect 6170 6614 6228 6624
rect 6556 7076 6614 7086
rect 6422 6626 6556 7058
rect 6364 6614 6422 6624
rect 6614 6814 6624 7058
rect 7074 6844 7196 7104
rect 7756 7104 7776 7282
rect 8020 7384 8872 7392
rect 8020 7378 9442 7384
rect 8020 7286 8408 7378
rect 7926 7270 8020 7280
rect 8464 7376 9442 7378
rect 8464 7286 8600 7376
rect 8408 7262 8464 7272
rect 8656 7374 9442 7376
rect 8656 7286 8802 7374
rect 8600 7260 8656 7270
rect 8858 7346 9442 7374
rect 8858 7268 9266 7346
rect 8802 7264 9266 7268
rect 8802 7258 8858 7264
rect 9244 7244 9266 7264
rect 9412 7340 9442 7346
rect 9412 7244 9440 7340
rect 10876 7336 10990 7342
rect 10872 7332 10990 7336
rect 10872 7326 10876 7332
rect 9244 7208 9440 7244
rect 9960 7276 10044 7286
rect 9244 7180 9442 7208
rect 10872 7238 10876 7242
rect 10872 7232 10990 7238
rect 10876 7228 10990 7232
rect 9960 7176 10044 7186
rect 8892 7152 8956 7158
rect 8512 7148 8956 7152
rect 8062 7144 8152 7148
rect 8058 7138 8152 7144
rect 8058 7134 8062 7138
rect 7756 7094 7764 7104
rect 7574 7064 7756 7074
rect 8512 7142 8892 7148
rect 8512 7140 8702 7142
rect 8512 7034 8514 7140
rect 8570 7036 8702 7140
rect 8758 7036 8892 7142
rect 8570 7034 8892 7036
rect 8512 7028 8892 7034
rect 8514 7012 8574 7028
rect 8702 7026 8758 7028
rect 10910 7100 10970 7108
rect 10592 7098 10972 7100
rect 8956 7028 8964 7070
rect 10592 7030 10910 7098
rect 10970 7030 10972 7098
rect 10592 7028 10972 7030
rect 8956 7024 8962 7028
rect 8892 7022 8962 7024
rect 8892 7014 8956 7022
rect 8058 6968 8062 6976
rect 8058 6966 8152 6968
rect 8062 6958 8152 6966
rect 10594 6998 10676 7028
rect 10910 7020 10970 7028
rect 7074 6814 7194 6844
rect 6614 6684 7196 6814
rect 7970 6792 8114 6802
rect 7970 6704 8114 6714
rect 9952 6724 10044 6734
rect 6614 6626 6624 6684
rect 6556 6610 6614 6620
rect 4626 6488 4902 6498
rect 4626 6044 4902 6054
rect 5882 5976 5940 5986
rect 5688 5966 5746 5976
rect 5654 5934 5688 5948
rect 5332 5842 5688 5934
rect 5746 5842 5882 5948
rect 5332 5642 5466 5842
rect 5532 5650 5882 5842
rect 5532 5642 5688 5650
rect 5332 5632 5688 5642
rect 5654 5514 5688 5632
rect 5746 5520 5882 5650
rect 6074 5974 6132 5984
rect 5940 5520 6074 5948
rect 5746 5518 6074 5520
rect 6266 5960 6324 5970
rect 6132 5518 6266 5948
rect 5746 5514 6266 5518
rect 5882 5510 5940 5514
rect 5688 5500 5746 5510
rect 6074 5508 6132 5514
rect 6458 5960 6516 5970
rect 6324 5514 6458 5948
rect 6266 5494 6324 5504
rect 6516 5514 6540 5948
rect 6458 5494 6516 5504
rect 4144 5124 4316 5126
rect 4142 5116 4232 5124
rect 4306 5116 4326 5124
rect 4142 4978 4144 5116
rect 4316 4978 4326 5116
rect 4142 4974 4326 4978
rect 7074 4986 7194 6684
rect 9952 6650 10044 6660
rect 10344 6548 10482 6558
rect 10344 6470 10482 6480
rect 8288 6382 8342 6392
rect 8276 6276 8288 6362
rect 8480 6382 8534 6392
rect 8342 6334 8480 6362
rect 8684 6362 8760 6364
rect 8534 6354 8770 6362
rect 8534 6334 8684 6354
rect 8342 6276 8476 6334
rect 8536 6282 8684 6334
rect 8760 6282 8770 6354
rect 8536 6276 8770 6282
rect 8476 6266 8480 6276
rect 8288 6246 8342 6256
rect 8534 6266 8536 6276
rect 8684 6272 8760 6276
rect 8480 6246 8534 6256
rect 7794 6234 7872 6244
rect 7794 6156 7872 6166
rect 10594 6150 10642 6998
rect 10866 6790 10996 6800
rect 10864 6778 10866 6788
rect 10988 6680 10996 6686
rect 10864 6676 10996 6680
rect 10864 6670 10988 6676
rect 7512 6134 7578 6144
rect 8178 6142 8244 6144
rect 8572 6142 8638 6144
rect 10594 6142 10678 6150
rect 8178 6134 8654 6142
rect 10100 6140 12748 6142
rect 10100 6136 10594 6140
rect 7578 6058 8178 6120
rect 8244 6132 8572 6134
rect 8244 6058 8376 6132
rect 7512 6056 8376 6058
rect 8442 6058 8572 6132
rect 8638 6058 8654 6134
rect 10072 6126 10594 6136
rect 9884 6120 10072 6122
rect 9874 6118 10072 6120
rect 8442 6056 8654 6058
rect 7512 6042 8654 6056
rect 9378 6062 9444 6072
rect 7512 6040 8244 6042
rect 7578 6020 8178 6040
rect 8376 6038 8442 6042
rect 8572 6040 8638 6042
rect 9378 5998 9380 6000
rect 9438 5998 9444 6000
rect 9378 5990 9444 5998
rect 9380 5988 9438 5990
rect 9114 5932 9166 5942
rect 9868 5930 10072 6118
rect 9166 5882 10072 5930
rect 10162 5888 10594 6126
rect 10678 6130 12748 6140
rect 10678 6124 12652 6130
rect 10678 5888 11110 6124
rect 10162 5882 11110 5888
rect 9166 5880 11110 5882
rect 9868 5878 11110 5880
rect 9868 5876 10226 5878
rect 9884 5874 10226 5876
rect 10072 5872 10162 5874
rect 11194 6116 12652 6124
rect 11194 5878 11628 6116
rect 9114 5858 9166 5868
rect 11110 5862 11194 5872
rect 11712 5878 12140 6116
rect 11628 5854 11712 5864
rect 12224 5878 12652 6116
rect 12736 5878 12748 6130
rect 12652 5868 12736 5878
rect 12140 5854 12224 5864
rect 9024 5726 9202 5736
rect 9024 5652 9202 5662
rect 7904 5398 8122 5408
rect 7904 5182 8122 5192
rect 10332 5134 10408 5188
rect 10846 5142 10950 5152
rect 10270 5122 10846 5134
rect 4144 4968 4316 4974
rect 6034 4878 6098 4888
rect 6034 4792 6098 4802
rect 6146 4868 6216 4878
rect 6204 4806 6216 4808
rect 6146 4798 6216 4806
rect 6146 4796 6204 4798
rect 7074 4760 7218 4986
rect 10246 4930 10340 5122
rect 10270 4924 10340 4930
rect 10416 4932 10846 5122
rect 11874 5138 11978 5148
rect 11370 5134 11474 5138
rect 10950 5128 11874 5134
rect 10950 4932 11370 5128
rect 10416 4924 11370 4932
rect 10270 4920 11370 4924
rect 10340 4914 10416 4920
rect 11474 4928 11874 5128
rect 12392 5142 12496 5152
rect 12290 5134 12392 5136
rect 11978 4932 12392 5134
rect 12496 5134 12600 5136
rect 12496 4932 12604 5134
rect 11978 4928 12604 4932
rect 11474 4920 12604 4928
rect 11874 4918 11978 4920
rect 11370 4908 11474 4918
rect 12290 4878 12600 4920
rect 5922 4740 7218 4760
rect 5922 4684 5926 4740
rect 5984 4684 7218 4740
rect 5922 4678 7218 4684
rect 5922 4672 7210 4678
rect 4230 4552 4304 4562
rect 4230 4464 4304 4474
<< via2 >>
rect 6782 10722 6998 10936
rect 4858 9944 5096 10320
rect 6558 10126 6560 10290
rect 6560 10126 6614 10290
rect 6614 10126 6628 10290
rect 6682 10262 6752 10282
rect 6682 10120 6732 10262
rect 6732 10120 6752 10262
rect 6682 10118 6752 10120
rect 11622 9866 11874 9868
rect 8946 9078 9022 9088
rect 8096 8966 8172 9002
rect 8096 8872 8098 8966
rect 8098 8872 8154 8966
rect 8154 8872 8172 8966
rect 8096 8860 8172 8872
rect 8946 8922 8958 9078
rect 8958 8922 9010 9078
rect 9010 8922 9022 9078
rect 8946 8918 9022 8922
rect 10356 9560 10424 9660
rect 11622 9454 11626 9866
rect 11626 9454 11874 9866
rect 9838 9436 9912 9450
rect 9838 9332 9848 9436
rect 9848 9332 9902 9436
rect 9902 9332 9912 9436
rect 9838 9324 9912 9332
rect 11606 8812 11888 9218
rect 7878 8178 7948 8286
rect 14292 7822 14338 7914
rect 14338 7822 14352 7914
rect 10876 7326 10990 7332
rect 9960 7186 10044 7276
rect 10876 7242 10970 7326
rect 10970 7242 10990 7326
rect 10876 7238 10990 7242
rect 8062 7134 8152 7138
rect 8062 6976 8152 7134
rect 8892 7024 8956 7148
rect 8062 6968 8152 6976
rect 4144 5024 4232 5116
rect 4232 5024 4306 5116
rect 4306 5024 4316 5116
rect 4144 4978 4316 5024
rect 9952 6660 10044 6724
rect 10344 6480 10482 6548
rect 8476 6276 8480 6334
rect 8480 6276 8534 6334
rect 8534 6276 8536 6334
rect 7806 6166 7860 6234
rect 7860 6166 7872 6234
rect 10864 6686 10866 6778
rect 10866 6686 10988 6778
rect 10864 6680 10988 6686
rect 9380 6000 9438 6054
rect 9380 5998 9438 6000
rect 9024 5662 9202 5726
rect 7904 5192 8122 5398
rect 6034 4860 6098 4878
rect 6034 4804 6092 4860
rect 6092 4804 6098 4860
rect 6034 4802 6098 4804
rect 6146 4862 6216 4868
rect 6146 4808 6204 4862
rect 6204 4808 6216 4862
rect 10340 4924 10416 5122
rect 4234 4480 4304 4550
<< metal3 >>
rect 6772 10936 7008 10941
rect 6772 10722 6782 10936
rect 6998 10722 7008 10936
rect 6772 10717 7008 10722
rect 4848 10320 5106 10325
rect 4848 9944 4858 10320
rect 5096 9944 5106 10320
rect 6548 10294 6638 10295
rect 6548 10290 6750 10294
rect 6548 10126 6558 10290
rect 6628 10287 6750 10290
rect 6628 10282 6762 10287
rect 6628 10126 6682 10282
rect 6548 10121 6682 10126
rect 6558 10118 6682 10121
rect 6752 10118 6762 10282
rect 6558 10113 6762 10118
rect 6558 10106 6750 10113
rect 4848 9939 5106 9944
rect 11612 9868 11884 9873
rect 10346 9660 10434 9665
rect 10346 9560 10356 9660
rect 10424 9560 10434 9660
rect 10346 9555 10434 9560
rect 9828 9450 9922 9455
rect 9828 9324 9838 9450
rect 9912 9324 9922 9450
rect 11612 9454 11622 9868
rect 11874 9454 11884 9868
rect 11612 9449 11884 9454
rect 9828 9319 9922 9324
rect 11606 9223 11910 9228
rect 11596 9218 11910 9223
rect 8936 9088 9032 9093
rect 8090 9007 8184 9020
rect 8086 9002 8184 9007
rect 8086 8860 8096 9002
rect 8172 8860 8184 9002
rect 8936 8918 8946 9088
rect 9022 8918 9032 9088
rect 8936 8913 9032 8918
rect 8086 8855 8184 8860
rect 8090 8676 8184 8855
rect 11596 8812 11606 9218
rect 11888 8812 11910 9218
rect 11596 8807 11910 8812
rect 11606 8676 11910 8807
rect 8088 8622 11948 8676
rect 8088 8566 9036 8622
rect 9130 8566 11948 8622
rect 8088 8476 11948 8566
rect 7050 8324 7444 8436
rect 7050 8286 7968 8324
rect 7050 8178 7878 8286
rect 7948 8178 7968 8286
rect 7050 8128 7968 8178
rect 4134 5116 4326 5121
rect 4134 4978 4144 5116
rect 4316 4978 4326 5116
rect 4134 4973 4326 4978
rect 6024 4882 6108 4883
rect 7050 4882 7444 8128
rect 14282 7822 14292 7920
rect 14370 7822 14380 7920
rect 14282 7817 14362 7822
rect 10866 7332 11000 7337
rect 9950 7276 10054 7281
rect 8894 7168 9006 7206
rect 9950 7186 9960 7276
rect 10044 7186 10054 7276
rect 10866 7238 10876 7332
rect 10990 7238 11000 7332
rect 10866 7233 11000 7238
rect 9950 7181 10054 7186
rect 8884 7148 9006 7168
rect 8052 7138 8162 7143
rect 8052 6968 8062 7138
rect 8152 6968 8162 7138
rect 8052 6963 8162 6968
rect 8882 7024 8892 7148
rect 8956 7140 9006 7148
rect 8956 7066 8998 7140
rect 8956 7024 9004 7066
rect 8882 6976 9004 7024
rect 7792 6234 7914 6846
rect 7792 6166 7806 6234
rect 7872 6166 7914 6234
rect 7792 6144 7914 6166
rect 8464 6334 8556 6386
rect 8464 6276 8476 6334
rect 8536 6276 8556 6334
rect 7894 5398 8132 5403
rect 7894 5396 7904 5398
rect 7854 5192 7904 5396
rect 8122 5396 8132 5398
rect 8122 5354 8136 5396
rect 8464 5354 8556 6276
rect 8882 5732 8970 6976
rect 10856 6784 10988 6798
rect 10856 6783 11008 6784
rect 10854 6778 11008 6783
rect 9938 6736 10070 6760
rect 10854 6736 10864 6778
rect 9938 6724 10864 6736
rect 9938 6660 9952 6724
rect 10044 6680 10864 6724
rect 10988 6680 11008 6778
rect 10044 6676 11008 6680
rect 10044 6672 11004 6676
rect 10044 6660 10988 6672
rect 9942 6655 10988 6660
rect 9944 6654 10988 6655
rect 9958 6642 10984 6654
rect 10334 6548 10492 6553
rect 10334 6480 10344 6548
rect 10482 6480 10492 6548
rect 10334 6475 10492 6480
rect 9376 6059 9468 6062
rect 9370 6054 9468 6059
rect 9370 5998 9380 6054
rect 9438 5998 9468 6054
rect 9370 5993 9468 5998
rect 9376 5946 9468 5993
rect 8882 5731 9102 5732
rect 8882 5726 9212 5731
rect 8882 5662 9024 5726
rect 9202 5662 9212 5726
rect 8882 5657 9212 5662
rect 8882 5598 9162 5657
rect 8882 5354 8970 5598
rect 9400 5354 9468 5946
rect 8122 5334 9178 5354
rect 9340 5334 9486 5354
rect 8122 5204 9486 5334
rect 8122 5192 8136 5204
rect 7854 4882 8136 5192
rect 8882 5178 8970 5204
rect 9102 5200 9422 5204
rect 10332 5127 10408 5188
rect 10330 5122 10426 5127
rect 10330 4924 10340 5122
rect 10416 4924 10426 5122
rect 10330 4919 10426 4924
rect 6024 4878 8162 4882
rect 6024 4802 6034 4878
rect 6098 4868 8162 4878
rect 6098 4808 6146 4868
rect 6216 4808 8162 4868
rect 6098 4802 8162 4808
rect 6024 4797 6108 4802
rect 4198 4550 4314 4566
rect 4198 4480 4234 4550
rect 4304 4480 4314 4550
rect 4198 4444 4314 4480
rect 7050 4444 7444 4802
rect 7854 4444 8136 4802
rect 4178 4242 8142 4444
rect 4590 4240 5020 4242
rect 7050 4238 7444 4242
rect 7854 4220 8136 4242
<< via3 >>
rect 6782 10722 6998 10936
rect 4858 9944 5096 10320
rect 6558 10126 6628 10290
rect 6682 10118 6752 10282
rect 10356 9560 10424 9660
rect 9838 9324 9912 9450
rect 11622 9454 11874 9868
rect 4144 4978 4316 5116
rect 14292 7914 14370 7920
rect 14292 7822 14352 7914
rect 14352 7822 14370 7914
rect 9960 7186 10044 7276
rect 10876 7238 10990 7332
rect 8062 6968 8152 7138
rect 7806 6166 7872 6234
rect 10344 6480 10482 6548
rect 10340 4924 10416 5122
<< metal4 >>
rect 4818 10950 5116 10954
rect 4748 10948 6976 10950
rect 4132 10937 6976 10948
rect 4132 10936 6999 10937
rect 4132 10734 6782 10936
rect 4132 10720 5116 10734
rect 6781 10722 6782 10734
rect 6998 10892 6999 10936
rect 7084 10892 7316 10902
rect 9552 10892 9912 10900
rect 6998 10802 9912 10892
rect 6998 10742 9916 10802
rect 6998 10740 9654 10742
rect 6998 10738 7780 10740
rect 7908 10738 9654 10740
rect 6998 10722 6999 10738
rect 6781 10721 6999 10722
rect 4142 5117 4296 10720
rect 4818 10320 5116 10720
rect 4818 9944 4858 10320
rect 5096 9944 5116 10320
rect 7084 10294 7316 10738
rect 9846 10294 9916 10742
rect 10876 10294 10994 10316
rect 11812 10294 12210 10296
rect 14288 10294 14386 10308
rect 6554 10290 7328 10294
rect 6554 10126 6558 10290
rect 6628 10282 7328 10290
rect 6628 10126 6682 10282
rect 6554 10124 6682 10126
rect 6556 10118 6682 10124
rect 6752 10124 7328 10282
rect 9766 10176 14386 10294
rect 6752 10122 6792 10124
rect 6752 10118 6753 10122
rect 6556 10117 6753 10118
rect 6556 10114 6752 10117
rect 4818 9910 5116 9944
rect 7084 6848 7316 10124
rect 9854 9451 9932 10176
rect 10336 10128 10480 10176
rect 9837 9450 9932 9451
rect 9837 9324 9838 9450
rect 9912 9324 9932 9450
rect 9837 9323 9932 9324
rect 9854 7404 9932 9323
rect 9850 7282 9932 7404
rect 10340 9660 10478 10128
rect 10340 9560 10356 9660
rect 10424 9560 10478 9660
rect 9850 7280 10040 7282
rect 9850 7276 10052 7280
rect 9850 7196 9960 7276
rect 9926 7188 9960 7196
rect 9959 7186 9960 7188
rect 10044 7188 10052 7276
rect 10044 7186 10045 7188
rect 9959 7185 10045 7186
rect 8056 7139 8116 7156
rect 8056 7138 8153 7139
rect 8056 6968 8062 7138
rect 8152 6968 8153 7138
rect 8056 6967 8153 6968
rect 8056 6848 8116 6967
rect 7084 6696 8202 6848
rect 10340 6834 10478 9560
rect 10876 7333 10994 10176
rect 11606 10170 12210 10176
rect 11606 9868 11882 10170
rect 11606 9458 11622 9868
rect 11621 9454 11622 9458
rect 11874 9458 11882 9868
rect 11874 9454 11875 9458
rect 11621 9453 11875 9454
rect 14288 7920 14386 10176
rect 14288 7822 14292 7920
rect 14370 7822 14386 7920
rect 14288 7804 14386 7822
rect 10875 7332 10994 7333
rect 10875 7238 10876 7332
rect 10990 7248 10994 7332
rect 10990 7238 10991 7248
rect 10875 7237 10991 7238
rect 7084 6690 7316 6696
rect 7730 6682 7914 6696
rect 7792 6234 7914 6682
rect 10340 6656 10482 6834
rect 7792 6166 7806 6234
rect 7872 6166 7914 6234
rect 7792 6144 7914 6166
rect 10342 6549 10482 6656
rect 10342 6548 10483 6549
rect 10342 6480 10344 6548
rect 10482 6480 10483 6548
rect 10342 6479 10483 6480
rect 10342 5188 10482 6479
rect 10332 5122 10482 5188
rect 4142 5116 4317 5117
rect 4142 5002 4144 5116
rect 4143 4978 4144 5002
rect 4316 4978 4317 5116
rect 4143 4977 4317 4978
rect 10339 4924 10340 5122
rect 10416 4926 10482 5122
rect 10416 4924 10478 4926
rect 10339 4923 10417 4924
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1723031900
transform 1 0 6017 0 1 4772
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_U2JGXT  sky130_fd_pr__nfet_01v8_U2JGXT_0
timestamp 1723031900
transform 0 1 8396 -1 0 8206
box -226 -510 226 510
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_0
timestamp 1723031900
transform 1 0 11752 0 1 9335
box -307 -704 307 704
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_1
timestamp 1723031900
transform 1 0 4959 0 1 9804
box -307 -704 307 704
use sky130_fd_pr__res_xhigh_po_1p41_VHK7CU  sky130_fd_pr__res_xhigh_po_1p41_VHK7CU_2
timestamp 1723031900
transform 1 0 4759 0 1 6622
box -307 -704 307 704
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723031900
transform 1 0 4070 0 1 4524
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1723031900
transform 1 0 10226 0 1 6688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1723031900
transform 1 0 10800 0 1 6696
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723031900
transform 1 0 4228 0 1 4520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  x5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723031900
transform 1 0 10892 0 1 6696
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1723031900
transform 1 0 9958 0 1 6688
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_BBNS5R  XM3
timestamp 1723031900
transform 1 0 8889 0 1 9654
box -359 -1110 359 1110
use sky130_fd_pr__pfet_01v8_SKB8VM  XM4
timestamp 1723031900
transform 1 0 6100 0 1 7975
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_SKB8VM  XM5
timestamp 1723031900
transform -1 0 6076 0 -1 9087
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_SKB8VM  XM6
timestamp 1723031900
transform -1 0 6056 0 -1 10179
box -696 -419 696 419
use sky130_fd_pr__pfet_01v8_VC5S4W  XM7
timestamp 1723031900
transform -1 0 6103 0 -1 6283
box -647 -1019 647 1019
use sky130_fd_pr__nfet_01v8_69TQ3K  XM8
timestamp 1723031900
transform 1 0 9268 0 1 5966
box -296 -310 296 310
use sky130_fd_pr__pfet_01v8_UGNVTG  XM9
timestamp 1723031900
transform -1 0 7809 0 -1 9641
box -359 -1119 359 1119
use sky130_fd_pr__pfet_01v8_XGS3BL  XM10
timestamp 1723031900
transform 1 0 10019 0 1 9509
box -407 -419 407 419
use sky130_fd_pr__nfet_01v8_MSLS59  XM11
timestamp 1723031900
transform 1 0 8407 0 1 6088
box -359 -510 359 510
use sky130_fd_pr__pfet_01v8_3HMWVM  XM12
timestamp 1723031900
transform 1 0 7684 0 1 6149
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_PDPE9S  XM13
timestamp 1723031900
transform 1 0 11409 0 1 5529
box -1457 -1019 1457 1019
use sky130_fd_pr__nfet_01v8_SC2JGL  XM14
timestamp 1723031900
transform 1 0 8681 0 1 7192
box -407 -410 407 410
use sky130_fd_pr__pfet_01v8_XGSNAL  XM15
timestamp 1723031900
transform 1 0 8039 0 1 7241
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_KRS3CJ  XM16
timestamp 1723031900
transform 1 0 11784 0 1 7869
box -2696 -319 2696 319
<< labels >>
flabel metal1 7576 7088 7776 7288 0 FreeSans 256 0 0 0 Va
port 1 nsew
flabel metal1 4362 7526 4562 7726 0 FreeSans 256 0 0 0 PAD
port 2 nsew
flabel via1 6786 10732 6986 10932 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 11630 7092 11828 7286 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 9240 7180 9436 7380 0 FreeSans 256 0 0 0 Vb
port 3 nsew
flabel via1 7904 5192 8104 5392 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
