magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_p >>
rect -77 981 -19 987
rect 115 981 173 987
rect -77 947 -65 981
rect 115 947 127 981
rect -77 941 -19 947
rect 115 941 173 947
rect -173 -947 -115 -941
rect 19 -947 77 -941
rect -173 -981 -161 -947
rect 19 -981 31 -947
rect -173 -987 -115 -981
rect 19 -987 77 -981
<< nwell >>
rect -359 -1119 359 1119
<< pmos >>
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
<< pdiff >>
rect -221 888 -159 900
rect -221 -888 -209 888
rect -175 -888 -159 888
rect -221 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 221 900
rect 159 -888 175 888
rect 209 -888 221 888
rect 159 -900 221 -888
<< pdiffc >>
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
<< nsubdiff >>
rect -323 1049 -227 1083
rect 227 1049 323 1083
rect -323 987 -289 1049
rect 289 987 323 1049
rect -323 -1049 -289 -987
rect 289 -1049 323 -987
rect -323 -1083 -227 -1049
rect 227 -1083 323 -1049
<< nsubdiffcont >>
rect -227 1049 227 1083
rect -323 -987 -289 987
rect 289 -987 323 987
rect -227 -1083 227 -1049
<< poly >>
rect -81 981 -15 997
rect -81 947 -65 981
rect -31 947 -15 981
rect -81 931 -15 947
rect 111 981 177 997
rect 111 947 127 981
rect 161 947 177 981
rect 111 931 177 947
rect -159 900 -129 926
rect -63 900 -33 931
rect 33 900 63 926
rect 129 900 159 931
rect -159 -931 -129 -900
rect -63 -926 -33 -900
rect 33 -931 63 -900
rect 129 -926 159 -900
rect -177 -947 -111 -931
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect -177 -997 -111 -981
rect 15 -947 81 -931
rect 15 -981 31 -947
rect 65 -981 81 -947
rect 15 -997 81 -981
<< polycont >>
rect -65 947 -31 981
rect 127 947 161 981
rect -161 -981 -127 -947
rect 31 -981 65 -947
<< locali >>
rect -323 1049 -227 1083
rect 227 1049 323 1083
rect -323 987 -289 1049
rect 289 987 323 1049
rect -81 947 -65 981
rect -31 947 -15 981
rect 111 947 127 981
rect 161 947 177 981
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect -177 -981 -161 -947
rect -127 -981 -111 -947
rect 15 -981 31 -947
rect 65 -981 81 -947
rect -323 -1049 -289 -987
rect 289 -1049 323 -987
rect -323 -1083 -227 -1049
rect 227 -1083 323 -1049
<< viali >>
rect -65 947 -31 981
rect 127 947 161 981
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect -161 -981 -127 -947
rect 31 -981 65 -947
<< metal1 >>
rect -77 981 -19 987
rect -77 947 -65 981
rect -31 947 -19 981
rect -77 941 -19 947
rect 115 981 173 987
rect 115 947 127 981
rect 161 947 173 981
rect 115 941 173 947
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect -173 -947 -115 -941
rect -173 -981 -161 -947
rect -127 -981 -115 -947
rect -173 -987 -115 -981
rect 19 -947 77 -941
rect 19 -981 31 -947
rect 65 -981 77 -947
rect 19 -987 77 -981
<< properties >>
string FIXED_BBOX -306 -1066 306 1066
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 9.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
