magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_p >>
rect -77 372 -19 378
rect 115 372 173 378
rect -77 338 -65 372
rect 115 338 127 372
rect -77 332 -19 338
rect 115 332 173 338
rect -173 -338 -115 -332
rect 19 -338 77 -332
rect -173 -372 -161 -338
rect 19 -372 31 -338
rect -173 -378 -115 -372
rect 19 -378 77 -372
<< pwell >>
rect -359 -510 359 510
<< nmos >>
rect -159 -300 -129 300
rect -63 -300 -33 300
rect 33 -300 63 300
rect 129 -300 159 300
<< ndiff >>
rect -221 288 -159 300
rect -221 -288 -209 288
rect -175 -288 -159 288
rect -221 -300 -159 -288
rect -129 288 -63 300
rect -129 -288 -113 288
rect -79 -288 -63 288
rect -129 -300 -63 -288
rect -33 288 33 300
rect -33 -288 -17 288
rect 17 -288 33 288
rect -33 -300 33 -288
rect 63 288 129 300
rect 63 -288 79 288
rect 113 -288 129 288
rect 63 -300 129 -288
rect 159 288 221 300
rect 159 -288 175 288
rect 209 -288 221 288
rect 159 -300 221 -288
<< ndiffc >>
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
<< psubdiff >>
rect -323 440 -227 474
rect 227 440 323 474
rect -323 378 -289 440
rect 289 378 323 440
rect -323 -440 -289 -378
rect 289 -440 323 -378
rect -323 -474 -227 -440
rect 227 -474 323 -440
<< psubdiffcont >>
rect -227 440 227 474
rect -323 -378 -289 378
rect 289 -378 323 378
rect -227 -474 227 -440
<< poly >>
rect -81 372 -15 388
rect -81 338 -65 372
rect -31 338 -15 372
rect -159 300 -129 326
rect -81 322 -15 338
rect 111 372 177 388
rect 111 338 127 372
rect 161 338 177 372
rect -63 300 -33 322
rect 33 300 63 326
rect 111 322 177 338
rect 129 300 159 322
rect -159 -322 -129 -300
rect -177 -338 -111 -322
rect -63 -326 -33 -300
rect 33 -322 63 -300
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect -177 -388 -111 -372
rect 15 -338 81 -322
rect 129 -326 159 -300
rect 15 -372 31 -338
rect 65 -372 81 -338
rect 15 -388 81 -372
<< polycont >>
rect -65 338 -31 372
rect 127 338 161 372
rect -161 -372 -127 -338
rect 31 -372 65 -338
<< locali >>
rect -323 440 -227 474
rect 227 440 323 474
rect -323 378 -289 440
rect 289 378 323 440
rect -81 338 -65 372
rect -31 338 -15 372
rect 111 338 127 372
rect 161 338 177 372
rect -209 288 -175 304
rect -209 -304 -175 -288
rect -113 288 -79 304
rect -113 -304 -79 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 79 288 113 304
rect 79 -304 113 -288
rect 175 288 209 304
rect 175 -304 209 -288
rect -177 -372 -161 -338
rect -127 -372 -111 -338
rect 15 -372 31 -338
rect 65 -372 81 -338
rect -323 -440 -289 -378
rect 289 -440 323 -378
rect -323 -474 -227 -440
rect 227 -474 323 -440
<< viali >>
rect -65 338 -31 372
rect 127 338 161 372
rect -209 -288 -175 288
rect -113 -288 -79 288
rect -17 -288 17 288
rect 79 -288 113 288
rect 175 -288 209 288
rect -161 -372 -127 -338
rect 31 -372 65 -338
<< metal1 >>
rect -77 372 -19 378
rect -77 338 -65 372
rect -31 338 -19 372
rect -77 332 -19 338
rect 115 372 173 378
rect 115 338 127 372
rect 161 338 173 372
rect 115 332 173 338
rect -215 288 -169 300
rect -215 -288 -209 288
rect -175 -288 -169 288
rect -215 -300 -169 -288
rect -119 288 -73 300
rect -119 -288 -113 288
rect -79 -288 -73 288
rect -119 -300 -73 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 73 288 119 300
rect 73 -288 79 288
rect 113 -288 119 288
rect 73 -300 119 -288
rect 169 288 215 300
rect 169 -288 175 288
rect 209 -288 215 288
rect 169 -300 215 -288
rect -173 -338 -115 -332
rect -173 -372 -161 -338
rect -127 -372 -115 -338
rect -173 -378 -115 -372
rect 19 -338 77 -332
rect 19 -372 31 -338
rect 65 -372 77 -338
rect 19 -378 77 -372
<< properties >>
string FIXED_BBOX -306 -457 306 457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
