magic
tech sky130A
magscale 1 2
timestamp 1722957601
<< error_p >>
rect -77 881 -19 887
rect 115 881 173 887
rect -77 847 -65 881
rect 115 847 127 881
rect -77 841 -19 847
rect 115 841 173 847
rect -173 -847 -115 -841
rect 19 -847 77 -841
rect -173 -881 -161 -847
rect 19 -881 31 -847
rect -173 -887 -115 -881
rect 19 -887 77 -881
<< nwell >>
rect -359 -1019 359 1019
<< pmos >>
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
<< pdiff >>
rect -221 788 -159 800
rect -221 -788 -209 788
rect -175 -788 -159 788
rect -221 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 221 800
rect 159 -788 175 788
rect 209 -788 221 788
rect 159 -800 221 -788
<< pdiffc >>
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
<< nsubdiff >>
rect -323 949 -227 983
rect 227 949 323 983
rect -323 887 -289 949
rect 289 887 323 949
rect -323 -949 -289 -887
rect 289 -949 323 -887
rect -323 -983 -227 -949
rect 227 -983 323 -949
<< nsubdiffcont >>
rect -227 949 227 983
rect -323 -887 -289 887
rect 289 -887 323 887
rect -227 -983 227 -949
<< poly >>
rect -81 881 -15 897
rect -81 847 -65 881
rect -31 847 -15 881
rect -81 831 -15 847
rect 111 881 177 897
rect 111 847 127 881
rect 161 847 177 881
rect 111 831 177 847
rect -159 800 -129 826
rect -63 800 -33 831
rect 33 800 63 826
rect 129 800 159 831
rect -159 -831 -129 -800
rect -63 -826 -33 -800
rect 33 -831 63 -800
rect 129 -826 159 -800
rect -177 -847 -111 -831
rect -177 -881 -161 -847
rect -127 -881 -111 -847
rect -177 -897 -111 -881
rect 15 -847 81 -831
rect 15 -881 31 -847
rect 65 -881 81 -847
rect 15 -897 81 -881
<< polycont >>
rect -65 847 -31 881
rect 127 847 161 881
rect -161 -881 -127 -847
rect 31 -881 65 -847
<< locali >>
rect -323 949 -227 983
rect 227 949 323 983
rect -323 887 -289 949
rect 289 887 323 949
rect -81 847 -65 881
rect -31 847 -15 881
rect 111 847 127 881
rect 161 847 177 881
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect -177 -881 -161 -847
rect -127 -881 -111 -847
rect 15 -881 31 -847
rect 65 -881 81 -847
rect -323 -949 -289 -887
rect 289 -949 323 -887
rect -323 -983 -227 -949
rect 227 -983 323 -949
<< viali >>
rect -65 847 -31 881
rect 127 847 161 881
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect -161 -881 -127 -847
rect 31 -881 65 -847
<< metal1 >>
rect -77 881 -19 887
rect -77 847 -65 881
rect -31 847 -19 881
rect -77 841 -19 847
rect 115 881 173 887
rect 115 847 127 881
rect 161 847 173 881
rect 115 841 173 847
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect -173 -847 -115 -841
rect -173 -881 -161 -847
rect -127 -881 -115 -847
rect -173 -887 -115 -881
rect 19 -847 77 -841
rect 19 -881 31 -847
rect 65 -881 77 -847
rect 19 -887 77 -881
<< properties >>
string FIXED_BBOX -306 -966 306 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
