magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_p >>
rect -125 281 -67 287
rect 67 281 125 287
rect -125 247 -113 281
rect 67 247 79 281
rect -125 241 -67 247
rect 67 241 125 247
rect -221 -247 -163 -241
rect -29 -247 29 -241
rect 163 -247 221 -241
rect -221 -281 -209 -247
rect -29 -281 -17 -247
rect 163 -281 175 -247
rect -221 -287 -163 -281
rect -29 -287 29 -281
rect 163 -287 221 -281
<< nwell >>
rect -407 -419 407 419
<< pmos >>
rect -207 -200 -177 200
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
rect 177 -200 207 200
<< pdiff >>
rect -269 188 -207 200
rect -269 -188 -257 188
rect -223 -188 -207 188
rect -269 -200 -207 -188
rect -177 188 -111 200
rect -177 -188 -161 188
rect -127 -188 -111 188
rect -177 -200 -111 -188
rect -81 188 -15 200
rect -81 -188 -65 188
rect -31 -188 -15 188
rect -81 -200 -15 -188
rect 15 188 81 200
rect 15 -188 31 188
rect 65 -188 81 188
rect 15 -200 81 -188
rect 111 188 177 200
rect 111 -188 127 188
rect 161 -188 177 188
rect 111 -200 177 -188
rect 207 188 269 200
rect 207 -188 223 188
rect 257 -188 269 188
rect 207 -200 269 -188
<< pdiffc >>
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
<< nsubdiff >>
rect -371 349 -275 383
rect 275 349 371 383
rect -371 287 -337 349
rect 337 287 371 349
rect -371 -349 -337 -287
rect 337 -349 371 -287
rect -371 -383 -275 -349
rect 275 -383 371 -349
<< nsubdiffcont >>
rect -275 349 275 383
rect -371 -287 -337 287
rect 337 -287 371 287
rect -275 -383 275 -349
<< poly >>
rect -129 281 -63 297
rect -129 247 -113 281
rect -79 247 -63 281
rect -129 231 -63 247
rect 63 281 129 297
rect 63 247 79 281
rect 113 247 129 281
rect 63 231 129 247
rect -207 200 -177 226
rect -111 200 -81 231
rect -15 200 15 226
rect 81 200 111 231
rect 177 200 207 226
rect -207 -231 -177 -200
rect -111 -226 -81 -200
rect -15 -231 15 -200
rect 81 -226 111 -200
rect 177 -231 207 -200
rect -225 -247 -159 -231
rect -225 -281 -209 -247
rect -175 -281 -159 -247
rect -225 -297 -159 -281
rect -33 -247 33 -231
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect -33 -297 33 -281
rect 159 -247 225 -231
rect 159 -281 175 -247
rect 209 -281 225 -247
rect 159 -297 225 -281
<< polycont >>
rect -113 247 -79 281
rect 79 247 113 281
rect -209 -281 -175 -247
rect -17 -281 17 -247
rect 175 -281 209 -247
<< locali >>
rect -371 349 -275 383
rect 275 349 371 383
rect -371 287 -337 349
rect 337 287 371 349
rect -129 247 -113 281
rect -79 247 -63 281
rect 63 247 79 281
rect 113 247 129 281
rect -257 188 -223 204
rect -257 -204 -223 -188
rect -161 188 -127 204
rect -161 -204 -127 -188
rect -65 188 -31 204
rect -65 -204 -31 -188
rect 31 188 65 204
rect 31 -204 65 -188
rect 127 188 161 204
rect 127 -204 161 -188
rect 223 188 257 204
rect 223 -204 257 -188
rect -225 -281 -209 -247
rect -175 -281 -159 -247
rect -33 -281 -17 -247
rect 17 -281 33 -247
rect 159 -281 175 -247
rect 209 -281 225 -247
rect -371 -349 -337 -287
rect 337 -349 371 -287
rect -371 -383 -275 -349
rect 275 -383 371 -349
<< viali >>
rect -113 247 -79 281
rect 79 247 113 281
rect -257 -188 -223 188
rect -161 -188 -127 188
rect -65 -188 -31 188
rect 31 -188 65 188
rect 127 -188 161 188
rect 223 -188 257 188
rect -209 -281 -175 -247
rect -17 -281 17 -247
rect 175 -281 209 -247
<< metal1 >>
rect -125 281 -67 287
rect -125 247 -113 281
rect -79 247 -67 281
rect -125 241 -67 247
rect 67 281 125 287
rect 67 247 79 281
rect 113 247 125 281
rect 67 241 125 247
rect -263 188 -217 200
rect -263 -188 -257 188
rect -223 -188 -217 188
rect -263 -200 -217 -188
rect -167 188 -121 200
rect -167 -188 -161 188
rect -127 -188 -121 188
rect -167 -200 -121 -188
rect -71 188 -25 200
rect -71 -188 -65 188
rect -31 -188 -25 188
rect -71 -200 -25 -188
rect 25 188 71 200
rect 25 -188 31 188
rect 65 -188 71 188
rect 25 -200 71 -188
rect 121 188 167 200
rect 121 -188 127 188
rect 161 -188 167 188
rect 121 -200 167 -188
rect 217 188 263 200
rect 217 -188 223 188
rect 257 -188 263 188
rect 217 -200 263 -188
rect -221 -247 -163 -241
rect -221 -281 -209 -247
rect -175 -281 -163 -247
rect -221 -287 -163 -281
rect -29 -247 29 -241
rect -29 -281 -17 -247
rect 17 -281 29 -247
rect -29 -287 29 -281
rect 163 -247 221 -241
rect 163 -281 175 -247
rect 209 -281 221 -247
rect 163 -287 221 -281
<< properties >>
string FIXED_BBOX -354 -366 354 366
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.0 l 0.15 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
