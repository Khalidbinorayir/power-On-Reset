magic
tech sky130A
magscale 1 2
timestamp 1722957601
<< error_p >>
rect -77 872 -19 878
rect 115 872 173 878
rect -77 838 -65 872
rect 115 838 127 872
rect -77 832 -19 838
rect 115 832 173 838
rect -173 -838 -115 -832
rect 19 -838 77 -832
rect -173 -872 -161 -838
rect 19 -872 31 -838
rect -173 -878 -115 -872
rect 19 -878 77 -872
<< pwell >>
rect -359 -1010 359 1010
<< nmos >>
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
<< ndiff >>
rect -221 788 -159 800
rect -221 -788 -209 788
rect -175 -788 -159 788
rect -221 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 221 800
rect 159 -788 175 788
rect 209 -788 221 788
rect 159 -800 221 -788
<< ndiffc >>
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
<< psubdiff >>
rect -323 940 -227 974
rect 227 940 323 974
rect -323 878 -289 940
rect 289 878 323 940
rect -323 -940 -289 -878
rect 289 -940 323 -878
rect -323 -974 -227 -940
rect 227 -974 323 -940
<< psubdiffcont >>
rect -227 940 227 974
rect -323 -878 -289 878
rect 289 -878 323 878
rect -227 -974 227 -940
<< poly >>
rect -81 872 -15 888
rect -81 838 -65 872
rect -31 838 -15 872
rect -159 800 -129 826
rect -81 822 -15 838
rect 111 872 177 888
rect 111 838 127 872
rect 161 838 177 872
rect -63 800 -33 822
rect 33 800 63 826
rect 111 822 177 838
rect 129 800 159 822
rect -159 -822 -129 -800
rect -177 -838 -111 -822
rect -63 -826 -33 -800
rect 33 -822 63 -800
rect -177 -872 -161 -838
rect -127 -872 -111 -838
rect -177 -888 -111 -872
rect 15 -838 81 -822
rect 129 -826 159 -800
rect 15 -872 31 -838
rect 65 -872 81 -838
rect 15 -888 81 -872
<< polycont >>
rect -65 838 -31 872
rect 127 838 161 872
rect -161 -872 -127 -838
rect 31 -872 65 -838
<< locali >>
rect -323 940 -227 974
rect 227 940 323 974
rect -323 878 -289 940
rect 289 878 323 940
rect -81 838 -65 872
rect -31 838 -15 872
rect 111 838 127 872
rect 161 838 177 872
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect -177 -872 -161 -838
rect -127 -872 -111 -838
rect 15 -872 31 -838
rect 65 -872 81 -838
rect -323 -940 -289 -878
rect 289 -940 323 -878
rect -323 -974 -227 -940
rect 227 -974 323 -940
<< viali >>
rect -65 838 -31 872
rect 127 838 161 872
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect -161 -872 -127 -838
rect 31 -872 65 -838
<< metal1 >>
rect -77 872 -19 878
rect -77 838 -65 872
rect -31 838 -19 872
rect -77 832 -19 838
rect 115 872 173 878
rect 115 838 127 872
rect 161 838 173 872
rect 115 832 173 838
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect -173 -838 -115 -832
rect -173 -872 -161 -838
rect -127 -872 -115 -838
rect -173 -878 -115 -872
rect 19 -838 77 -832
rect 19 -872 31 -838
rect 65 -872 77 -838
rect 19 -878 77 -872
<< properties >>
string FIXED_BBOX -306 -957 306 957
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
