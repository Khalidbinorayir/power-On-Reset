* NGSPICE file created from por.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_VHK7CU a_n141_n538# a_n271_n668# a_n141_106#
X0 a_n141_106# a_n141_n538# a_n271_n668# sky130_fd_pr__res_xhigh_po_1p41 l=1.22
C0 a_n141_106# a_n141_n538# 0.073123f
C1 a_n141_n538# a_n271_n668# 0.770781f
C2 a_n141_106# a_n271_n668# 0.770781f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HMWVM w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ VSUBS
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 w_n296_n319# a_n158_n100# 0.085221f
C1 a_n158_n100# a_100_n100# 0.055609f
C2 a_n100_n197# a_n158_n100# 0.026809f
C3 w_n296_n319# a_100_n100# 0.085221f
C4 a_n100_n197# w_n296_n319# 0.434431f
C5 a_n100_n197# a_100_n100# 0.026809f
C6 a_100_n100# VSUBS 0.060699f
C7 a_n158_n100# VSUBS 0.060699f
C8 a_n100_n197# VSUBS 0.310981f
C9 w_n296_n319# VSUBS 1.64714f
.ends

.subckt sky130_fd_pr__pfet_01v8_PDPE9S a_1261_n800# a_29_n897# a_n1319_n800# a_n287_n800#
+ a_n745_n897# a_n1061_n800# a_745_n800# a_803_n897# a_n229_n897# a_n1003_n897# a_287_n897#
+ a_229_n800# w_n1457_n1019# a_n545_n800# a_1061_n897# a_1003_n800# a_n487_n897# a_n1261_n897#
+ a_n29_n800# a_487_n800# a_545_n897# a_n803_n800# VSUBS
X0 a_487_n800# a_287_n897# a_229_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X1 a_745_n800# a_545_n897# a_487_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2 a_1261_n800# a_1061_n897# a_1003_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X3 a_229_n800# a_29_n897# a_n29_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X4 a_n29_n800# a_n229_n897# a_n287_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X5 a_n545_n800# a_n745_n897# a_n803_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X6 a_n287_n800# a_n487_n897# a_n545_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X7 a_n803_n800# a_n1003_n897# a_n1061_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X8 a_n1061_n800# a_n1261_n897# a_n1319_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X9 a_1003_n800# a_803_n897# a_745_n800# w_n1457_n1019# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
C0 w_n1457_n1019# a_n29_n800# 0.021376f
C1 w_n1457_n1019# a_n287_n800# 0.021376f
C2 w_n1457_n1019# a_229_n800# 0.021376f
C3 a_487_n800# a_287_n897# 0.176406f
C4 a_n1261_n897# a_n1319_n800# 0.176406f
C5 a_29_n897# w_n1457_n1019# 0.353669f
C6 w_n1457_n1019# a_803_n897# 0.353893f
C7 a_1003_n800# a_745_n800# 0.437576f
C8 a_n487_n897# a_n287_n800# 0.176406f
C9 a_n803_n800# a_n545_n800# 0.437576f
C10 w_n1457_n1019# a_1003_n800# 0.021376f
C11 a_487_n800# a_545_n897# 0.176406f
C12 w_n1457_n1019# a_287_n897# 0.353666f
C13 a_n1003_n897# a_n803_n800# 0.176406f
C14 a_745_n800# a_545_n897# 0.176406f
C15 a_n1061_n800# a_n803_n800# 0.437576f
C16 w_n1457_n1019# a_n229_n897# 0.353669f
C17 a_n29_n800# a_n287_n800# 0.437576f
C18 a_n29_n800# a_229_n800# 0.437576f
C19 a_803_n897# a_1061_n897# 0.109462f
C20 w_n1457_n1019# a_n545_n800# 0.021376f
C21 a_487_n800# a_745_n800# 0.437576f
C22 a_n1003_n897# a_n1061_n800# 0.176406f
C23 w_n1457_n1019# a_545_n897# 0.353723f
C24 a_29_n897# a_n29_n800# 0.176406f
C25 a_n745_n897# a_n545_n800# 0.176406f
C26 a_29_n897# a_229_n800# 0.176406f
C27 a_1261_n800# w_n1457_n1019# 0.512046f
C28 a_n487_n897# a_n229_n897# 0.109462f
C29 w_n1457_n1019# a_n803_n800# 0.021376f
C30 a_487_n800# w_n1457_n1019# 0.021376f
C31 a_n745_n897# a_n803_n800# 0.176406f
C32 a_1003_n800# a_1061_n897# 0.176406f
C33 a_n487_n897# a_n545_n800# 0.176406f
C34 w_n1457_n1019# a_n1003_n897# 0.353893f
C35 w_n1457_n1019# a_n1061_n800# 0.021376f
C36 a_n1003_n897# a_n745_n897# 0.109462f
C37 w_n1457_n1019# a_745_n800# 0.021376f
C38 a_803_n897# a_1003_n800# 0.176406f
C39 a_287_n897# a_229_n800# 0.176406f
C40 a_n29_n800# a_n229_n897# 0.176406f
C41 a_n287_n800# a_n229_n897# 0.176406f
C42 a_29_n897# a_287_n897# 0.109462f
C43 a_n1261_n897# a_n1003_n897# 0.109462f
C44 a_n1261_n897# a_n1061_n800# 0.176406f
C45 w_n1457_n1019# a_n745_n897# 0.353723f
C46 a_29_n897# a_n229_n897# 0.109462f
C47 a_n287_n800# a_n545_n800# 0.437576f
C48 a_1261_n800# a_1061_n897# 0.176406f
C49 a_n1061_n800# a_n1319_n800# 0.437576f
C50 a_803_n897# a_545_n897# 0.109462f
C51 w_n1457_n1019# a_n487_n897# 0.353666f
C52 a_487_n800# a_229_n800# 0.437576f
C53 a_n1261_n897# w_n1457_n1019# 0.394013f
C54 a_n745_n897# a_n487_n897# 0.109462f
C55 w_n1457_n1019# a_n1319_n800# 0.512046f
C56 a_1261_n800# a_1003_n800# 0.437576f
C57 w_n1457_n1019# a_1061_n897# 0.394013f
C58 a_287_n897# a_545_n897# 0.109462f
C59 a_803_n897# a_745_n800# 0.176406f
C60 a_1261_n800# VSUBS 0.413693f
C61 a_1003_n800# VSUBS 0.227763f
C62 a_745_n800# VSUBS 0.227763f
C63 a_487_n800# VSUBS 0.227763f
C64 a_229_n800# VSUBS 0.227763f
C65 a_n29_n800# VSUBS 0.227763f
C66 a_n287_n800# VSUBS 0.227763f
C67 a_n545_n800# VSUBS 0.227763f
C68 a_n803_n800# VSUBS 0.227763f
C69 a_n1061_n800# VSUBS 0.227763f
C70 a_n1319_n800# VSUBS 0.413693f
C71 a_1061_n897# VSUBS 0.335881f
C72 a_803_n897# VSUBS 0.307579f
C73 a_545_n897# VSUBS 0.307579f
C74 a_287_n897# VSUBS 0.307579f
C75 a_29_n897# VSUBS 0.307579f
C76 a_n229_n897# VSUBS 0.307579f
C77 a_n487_n897# VSUBS 0.307579f
C78 a_n745_n897# VSUBS 0.307579f
C79 a_n1003_n897# VSUBS 0.307579f
C80 a_n1261_n897# VSUBS 0.335881f
C81 w_n1457_n1019# VSUBS 20.2216f
.ends

.subckt sky130_fd_pr__nfet_01v8_SC2JGL a_15_n200# a_n177_n200# a_111_n200# a_159_n288#
+ a_63_222# a_n81_n200# a_n129_222# a_n269_n200# a_207_n200# a_n225_n288# a_n371_n374#
+ a_n33_n288#
X0 a_n81_n200# a_n129_222# a_n177_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X1 a_15_n200# a_n33_n288# a_n81_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X2 a_207_n200# a_159_n288# a_111_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X3 a_n177_n200# a_n225_n288# a_n269_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X4 a_111_n200# a_63_222# a_15_n200# a_n371_n374# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
C0 a_159_n288# a_n33_n288# 0.02473f
C1 a_n269_n200# a_n177_n200# 0.296004f
C2 a_159_n288# a_111_n200# 0.017011f
C3 a_n81_n200# a_n129_222# 0.017011f
C4 a_63_222# a_15_n200# 0.017011f
C5 a_n129_222# a_n225_n288# 0.013333f
C6 a_111_n200# a_207_n200# 0.296004f
C7 a_63_222# a_n33_n288# 0.013333f
C8 a_15_n200# a_n33_n288# 0.017011f
C9 a_63_222# a_111_n200# 0.017011f
C10 a_15_n200# a_111_n200# 0.296004f
C11 a_n81_n200# a_n177_n200# 0.296004f
C12 a_n129_222# a_n177_n200# 0.017011f
C13 a_n225_n288# a_n177_n200# 0.017011f
C14 a_15_n200# a_n81_n200# 0.296004f
C15 a_n269_n200# a_n225_n288# 0.017011f
C16 a_63_222# a_n129_222# 0.02473f
C17 a_n81_n200# a_n33_n288# 0.017011f
C18 a_159_n288# a_207_n200# 0.017011f
C19 a_n129_222# a_n33_n288# 0.013333f
C20 a_n33_n288# a_n225_n288# 0.02473f
C21 a_63_222# a_159_n288# 0.013333f
C22 a_207_n200# a_n371_n374# 0.238762f
C23 a_111_n200# a_n371_n374# 0.047715f
C24 a_15_n200# a_n371_n374# 0.047715f
C25 a_n81_n200# a_n371_n374# 0.047715f
C26 a_n177_n200# a_n371_n374# 0.047715f
C27 a_n269_n200# a_n371_n374# 0.238762f
C28 a_159_n288# a_n371_n374# 0.184753f
C29 a_n33_n288# a_n371_n374# 0.153467f
C30 a_63_222# a_n371_n374# 0.172901f
C31 a_n225_n288# a_n371_n374# 0.184753f
C32 a_n129_222# a_n371_n374# 0.172901f
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 VGND A 0.040045f
C1 VPB Y 0.017744f
C2 VPB VPWR 0.054478f
C3 A Y 0.047605f
C4 A VPWR 0.037031f
C5 VPB A 0.045062f
C6 VGND Y 0.099841f
C7 VGND VPWR 0.033816f
C8 Y VPWR 0.127579f
C9 VGND VPB 0.009478f
C10 VGND VNB 0.251126f
C11 Y VNB 0.096099f
C12 VPWR VNB 0.218922f
C13 A VNB 0.166643f
C14 VPB VNB 0.338976f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGSNAL a_n33_n397# a_n73_n300# a_15_n300# w_n211_n519#
+ VSUBS
X0 a_15_n300# a_n33_n397# a_n73_n300# w_n211_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
C0 w_n211_n519# a_15_n300# 0.203636f
C1 w_n211_n519# a_n73_n300# 0.203636f
C2 a_n33_n397# a_15_n300# 0.034115f
C3 a_n33_n397# a_n73_n300# 0.034115f
C4 w_n211_n519# a_n33_n397# 0.241085f
C5 a_15_n300# a_n73_n300# 0.479983f
C6 a_15_n300# VSUBS 0.130707f
C7 a_n73_n300# VSUBS 0.130707f
C8 a_n33_n397# VSUBS 0.120511f
C9 w_n211_n519# VSUBS 1.93133f
.ends

.subckt sky130_fd_pr__nfet_01v8_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
C0 a_n33_n188# a_15_n100# 0.025448f
C1 a_n73_n100# a_15_n100# 0.162113f
C2 a_n33_n188# a_n73_n100# 0.025448f
C3 a_15_n100# a_n175_n274# 0.131704f
C4 a_n73_n100# a_n175_n274# 0.131704f
C5 a_n33_n188# a_n175_n274# 0.34289f
.ends

.subckt sky130_fd_pr__pfet_01v8_KRS3CJ a_n2500_n197# a_2500_n100# a_n2558_n100# w_n2696_n319#
+ VSUBS
X0 a_2500_n100# a_n2500_n197# a_n2558_n100# w_n2696_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=25
C0 w_n2696_n319# a_2500_n100# 0.085193f
C1 w_n2696_n319# a_n2558_n100# 0.085193f
C2 a_n2500_n197# a_2500_n100# 0.049339f
C3 a_n2500_n197# a_n2558_n100# 0.049339f
C4 w_n2696_n319# a_n2500_n197# 7.83378f
C5 a_2500_n100# VSUBS 0.091337f
C6 a_n2558_n100# VSUBS 0.091337f
C7 a_n2500_n197# VSUBS 6.64706f
C8 w_n2696_n319# VSUBS 13.1108f
.ends

.subckt sky130_fd_sc_hd__and2_0 A B VGND VNB VPB VPWR X a_123_47# a_40_47#
X0 VPWR B a_40_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1841 pd=1.26 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_40_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1696 pd=1.81 as=0.1841 ps=1.26 w=0.64 l=0.15
X2 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0966 pd=0.88 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 X a_40_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0966 ps=0.88 w=0.42 l=0.15
X4 a_123_47# A a_40_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1113 ps=1.37 w=0.42 l=0.15
X5 a_40_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1113 ps=1.37 w=0.42 l=0.15
C0 VPB X 0.022086f
C1 A VPWR 0.047791f
C2 VPB VPWR 0.062434f
C3 VPWR X 0.111278f
C4 a_40_47# VGND 0.138964f
C5 a_123_47# X 2.99e-19
C6 a_123_47# VPWR 5.63e-19
C7 B a_40_47# 0.206108f
C8 B VGND 0.019565f
C9 a_40_47# A 0.12536f
C10 a_40_47# VPB 0.082909f
C11 VGND A 0.017409f
C12 a_40_47# X 0.11426f
C13 VGND VPB 0.006814f
C14 B A 0.117044f
C15 a_40_47# VPWR 0.141098f
C16 B VPB 0.088046f
C17 VGND X 0.105358f
C18 a_123_47# a_40_47# 0.004822f
C19 VGND VPWR 0.045704f
C20 B X 0.007578f
C21 B VPWR 0.044651f
C22 a_123_47# VGND 0.00394f
C23 A VPB 0.093286f
C24 A X 1.67e-19
C25 VGND VNB 0.300193f
C26 X VNB 0.10272f
C27 VPWR VNB 0.262881f
C28 B VNB 0.121465f
C29 A VNB 0.194569f
C30 VPB VNB 0.516168f
C31 a_40_47# VNB 0.230074f
.ends

.subckt sky130_fd_pr__nfet_01v8_BBNS5R a_n33_n900# a_15_n988# a_n81_922# a_n177_n988#
+ a_159_n900# a_n221_n900# a_n129_n900# a_63_n900# a_111_922# a_n323_n1074#
X0 a_n33_n900# a_n81_922# a_n129_n900# a_n323_n1074# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X1 a_159_n900# a_111_922# a_63_n900# a_n323_n1074# sky130_fd_pr__nfet_01v8 ad=2.79 pd=18.62 as=1.485 ps=9.33 w=9 l=0.15
X2 a_63_n900# a_15_n988# a_n33_n900# a_n323_n1074# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X3 a_n129_n900# a_n177_n988# a_n221_n900# a_n323_n1074# sky130_fd_pr__nfet_01v8 ad=1.485 pd=9.33 as=2.79 ps=18.62 w=9 l=0.15
C0 a_n129_n900# a_n33_n900# 1.32129f
C1 a_111_922# a_159_n900# 0.045972f
C2 a_15_n988# a_n33_n900# 0.045972f
C3 a_n81_922# a_n177_n988# 0.013333f
C4 a_111_922# a_15_n988# 0.013333f
C5 a_n221_n900# a_n177_n988# 0.045972f
C6 a_63_n900# a_n33_n900# 1.32129f
C7 a_111_922# a_63_n900# 0.045972f
C8 a_n129_n900# a_n81_922# 0.045972f
C9 a_159_n900# a_63_n900# 1.32129f
C10 a_n129_n900# a_n177_n988# 0.045972f
C11 a_n81_922# a_n33_n900# 0.045972f
C12 a_111_922# a_n81_922# 0.02473f
C13 a_63_n900# a_15_n988# 0.045972f
C14 a_15_n988# a_n81_922# 0.013333f
C15 a_n129_n900# a_n221_n900# 1.32129f
C16 a_15_n988# a_n177_n988# 0.02473f
C17 a_159_n900# a_n323_n1074# 0.952557f
C18 a_63_n900# a_n323_n1074# 0.106844f
C19 a_n33_n900# a_n323_n1074# 0.106844f
C20 a_n129_n900# a_n323_n1074# 0.106844f
C21 a_n221_n900# a_n323_n1074# 0.952557f
C22 a_15_n988# a_n323_n1074# 0.170096f
C23 a_111_922# a_n323_n1074# 0.181931f
C24 a_n177_n988# a_n323_n1074# 0.181931f
C25 a_n81_922# a_n323_n1074# 0.170096f
.ends

.subckt sky130_fd_pr__pfet_01v8_SKB8VM w_n696_n419# a_n500_n297# a_500_n200# a_n558_n200#
+ VSUBS
X0 a_500_n200# a_n500_n297# a_n558_n200# w_n696_n419# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=5
C0 a_n500_n297# a_500_n200# 0.086192f
C1 a_n558_n200# a_500_n200# 0.026656f
C2 w_n696_n419# a_500_n200# 0.146171f
C3 a_n500_n297# a_n558_n200# 0.086192f
C4 a_n500_n297# w_n696_n419# 1.66884f
C5 w_n696_n419# a_n558_n200# 0.146171f
C6 a_500_n200# VSUBS 0.144387f
C7 a_n558_n200# VSUBS 0.144387f
C8 a_n500_n297# VSUBS 1.43114f
C9 w_n696_n419# VSUBS 4.49444f
.ends

.subckt sky130_fd_pr__pfet_01v8_VC5S4W w_n647_n1019# a_63_n800# a_n225_n800# a_399_831#
+ a_111_n897# a_n321_n800# a_n273_n897# a_15_831# a_207_831# a_n33_n800# a_n509_n800#
+ a_447_n800# a_n81_n897# a_n177_831# a_159_n800# a_255_n800# a_n369_831# a_351_n800#
+ a_n417_n800# a_303_n897# a_n129_n800# a_n465_n897# VSUBS
X0 a_n33_n800# a_n81_n897# a_n129_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X1 a_351_n800# a_303_n897# a_255_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X2 a_255_n800# a_207_831# a_159_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X3 a_n321_n800# a_n369_831# a_n417_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X4 a_159_n800# a_111_n897# a_63_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X5 a_n225_n800# a_n273_n897# a_n321_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X6 a_447_n800# a_399_831# a_351_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=2.48 pd=16.62 as=1.32 ps=8.33 w=8 l=0.15
X7 a_63_n800# a_15_831# a_n33_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X8 a_n129_n800# a_n177_831# a_n225_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.15
X9 a_n417_n800# a_n465_n897# a_n509_n800# w_n647_n1019# sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=2.48 ps=16.62 w=8 l=0.15
C0 a_447_n800# w_n647_n1019# 0.51136f
C1 w_n647_n1019# a_n129_n800# 0.020004f
C2 a_n129_n800# a_n225_n800# 1.17482f
C3 a_n369_831# a_n321_n800# 0.041475f
C4 a_n417_n800# a_n369_831# 0.041475f
C5 a_n177_831# a_n81_n897# 0.012606f
C6 a_303_n897# a_207_831# 0.012606f
C7 a_n417_n800# a_n509_n800# 1.17482f
C8 a_n465_n897# a_n273_n897# 0.025732f
C9 w_n647_n1019# a_n225_n800# 0.020004f
C10 a_n129_n800# a_n81_n897# 0.041475f
C11 a_399_831# a_351_n800# 0.041475f
C12 a_255_n800# a_207_831# 0.041475f
C13 a_399_831# a_447_n800# 0.041475f
C14 w_n647_n1019# a_63_n800# 0.020004f
C15 a_255_n800# a_159_n800# 1.17482f
C16 w_n647_n1019# a_n81_n897# 0.108905f
C17 a_n369_831# a_n273_n897# 0.012606f
C18 w_n647_n1019# a_111_n897# 0.108917f
C19 a_n465_n897# a_n369_831# 0.012606f
C20 a_399_831# w_n647_n1019# 0.12444f
C21 a_n465_n897# a_n509_n800# 0.041475f
C22 a_63_n800# a_111_n897# 0.041475f
C23 a_n177_831# a_15_831# 0.025732f
C24 a_n81_n897# a_111_n897# 0.025732f
C25 a_303_n897# a_255_n800# 0.041475f
C26 w_n647_n1019# a_n321_n800# 0.020004f
C27 a_n321_n800# a_n225_n800# 1.17482f
C28 a_n417_n800# w_n647_n1019# 0.020004f
C29 a_n177_831# a_n273_n897# 0.012606f
C30 a_n129_n800# a_n33_n800# 1.17482f
C31 w_n647_n1019# a_207_831# 0.108947f
C32 w_n647_n1019# a_n33_n800# 0.020004f
C33 w_n647_n1019# a_159_n800# 0.020004f
C34 w_n647_n1019# a_15_831# 0.108905f
C35 a_303_n897# a_351_n800# 0.041475f
C36 a_n369_831# a_n177_831# 0.025732f
C37 a_n33_n800# a_63_n800# 1.17482f
C38 a_207_831# a_111_n897# 0.012606f
C39 w_n647_n1019# a_n273_n897# 0.108947f
C40 a_n225_n800# a_n273_n897# 0.041475f
C41 a_159_n800# a_63_n800# 1.17482f
C42 a_63_n800# a_15_831# 0.041475f
C43 a_n33_n800# a_n81_n897# 0.041475f
C44 a_n465_n897# w_n647_n1019# 0.12444f
C45 a_n81_n897# a_15_831# 0.012606f
C46 a_159_n800# a_111_n897# 0.041475f
C47 a_15_831# a_111_n897# 0.012606f
C48 a_399_831# a_207_831# 0.025732f
C49 a_255_n800# a_351_n800# 1.17482f
C50 a_n417_n800# a_n321_n800# 1.17482f
C51 a_303_n897# w_n647_n1019# 0.119704f
C52 a_n81_n897# a_n273_n897# 0.025732f
C53 a_n369_831# w_n647_n1019# 0.119704f
C54 w_n647_n1019# a_n509_n800# 0.51136f
C55 a_255_n800# w_n647_n1019# 0.020004f
C56 a_303_n897# a_111_n897# 0.025732f
C57 a_n129_n800# a_n177_831# 0.041475f
C58 a_447_n800# a_351_n800# 1.17482f
C59 a_303_n897# a_399_831# 0.012606f
C60 a_n321_n800# a_n273_n897# 0.041475f
C61 a_159_n800# a_207_831# 0.041475f
C62 a_207_831# a_15_831# 0.025732f
C63 a_n33_n800# a_15_831# 0.041475f
C64 a_n465_n897# a_n417_n800# 0.041475f
C65 w_n647_n1019# a_n177_831# 0.108917f
C66 a_n177_831# a_n225_n800# 0.041475f
C67 w_n647_n1019# a_351_n800# 0.020004f
C68 a_447_n800# VSUBS 0.338824f
C69 a_351_n800# VSUBS 0.078026f
C70 a_255_n800# VSUBS 0.078026f
C71 a_159_n800# VSUBS 0.078026f
C72 a_63_n800# VSUBS 0.078026f
C73 a_n33_n800# VSUBS 0.078026f
C74 a_n129_n800# VSUBS 0.078026f
C75 a_n225_n800# VSUBS 0.078026f
C76 a_n321_n800# VSUBS 0.078026f
C77 a_n417_n800# VSUBS 0.078026f
C78 a_n509_n800# VSUBS 0.338824f
C79 a_303_n897# VSUBS 0.055715f
C80 a_111_n897# VSUBS 0.046052f
C81 a_n81_n897# VSUBS 0.046052f
C82 a_n273_n897# VSUBS 0.046052f
C83 a_n465_n897# VSUBS 0.06269f
C84 a_399_831# VSUBS 0.06269f
C85 a_207_831# VSUBS 0.046052f
C86 a_15_831# VSUBS 0.046052f
C87 a_n177_831# VSUBS 0.046052f
C88 a_n369_831# VSUBS 0.055715f
C89 w_n647_n1019# VSUBS 9.5697f
.ends

.subckt sky130_fd_pr__nfet_01v8_69TQ3K a_n260_n274# a_100_n100# a_n158_n100# a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n260_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n188# a_n158_n100# 0.026809f
C1 a_100_n100# a_n158_n100# 0.055609f
C2 a_100_n100# a_n100_n188# 0.026809f
C3 a_100_n100# a_n260_n274# 0.146358f
C4 a_n158_n100# a_n260_n274# 0.146358f
C5 a_n100_n188# a_n260_n274# 0.724275f
.ends

.subckt sky130_fd_pr__pfet_01v8_UGNVTG a_n33_n900# a_159_n900# a_111_931# a_n221_n900#
+ a_n129_n900# w_n359_n1119# a_63_n900# a_15_n997# a_n81_931# a_n177_n997# VSUBS
X0 a_159_n900# a_111_931# a_63_n900# w_n359_n1119# sky130_fd_pr__pfet_01v8 ad=2.79 pd=18.62 as=1.485 ps=9.33 w=9 l=0.15
X1 a_63_n900# a_15_n997# a_n33_n900# w_n359_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
X2 a_n129_n900# a_n177_n997# a_n221_n900# w_n359_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=2.79 ps=18.62 w=9 l=0.15
X3 a_n33_n900# a_n81_931# a_n129_n900# w_n359_n1119# sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.15
C0 w_n359_n1119# a_n33_n900# 0.020004f
C1 a_n221_n900# a_n129_n900# 1.32129f
C2 a_n81_931# a_15_n997# 0.012606f
C3 a_63_n900# a_15_n997# 0.045418f
C4 a_n177_n997# w_n359_n1119# 0.124487f
C5 a_n81_931# a_n129_n900# 0.045418f
C6 a_63_n900# a_159_n900# 1.32129f
C7 w_n359_n1119# a_15_n997# 0.119783f
C8 a_n221_n900# w_n359_n1119# 0.572335f
C9 a_111_931# a_15_n997# 0.012606f
C10 a_15_n997# a_n33_n900# 0.045418f
C11 w_n359_n1119# a_n129_n900# 0.020004f
C12 w_n359_n1119# a_n81_931# 0.119783f
C13 a_n129_n900# a_n33_n900# 1.32129f
C14 a_111_931# a_n81_931# 0.025732f
C15 w_n359_n1119# a_63_n900# 0.020004f
C16 w_n359_n1119# a_159_n900# 0.572335f
C17 a_111_931# a_63_n900# 0.045418f
C18 a_111_931# a_159_n900# 0.045418f
C19 a_n177_n997# a_15_n997# 0.025732f
C20 a_n221_n900# a_n177_n997# 0.045418f
C21 a_n81_931# a_n33_n900# 0.045418f
C22 a_63_n900# a_n33_n900# 1.32129f
C23 a_n177_n997# a_n129_n900# 0.045418f
C24 a_n177_n997# a_n81_931# 0.012606f
C25 a_111_931# w_n359_n1119# 0.124487f
C26 a_159_n900# VSUBS 0.37982f
C27 a_63_n900# VSUBS 0.086473f
C28 a_n33_n900# VSUBS 0.086473f
C29 a_n129_n900# VSUBS 0.086473f
C30 a_n221_n900# VSUBS 0.37982f
C31 a_15_n997# VSUBS 0.055715f
C32 a_n177_n997# VSUBS 0.06269f
C33 a_111_931# VSUBS 0.06269f
C34 a_n81_931# VSUBS 0.055715f
C35 w_n359_n1119# VSUBS 6.22307f
.ends

.subckt sky130_fd_pr__nfet_01v8_U2JGXT a_30_n300# a_n88_n300# a_n33_n388# a_n190_n474#
X0 a_30_n300# a_n33_n388# a_n88_n300# a_n190_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.3
C0 a_n33_n388# a_n88_n300# 0.02692f
C1 a_30_n300# a_n33_n388# 0.02692f
C2 a_30_n300# a_n88_n300# 0.358546f
C3 a_30_n300# a_n190_n474# 0.346088f
C4 a_n88_n300# a_n190_n474# 0.346088f
C5 a_n33_n388# a_n190_n474# 0.350472f
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_15_n200# a_n177_n200# a_n129_231# a_111_n200#
+ w_n407_n419# a_n225_n297# a_n81_n200# a_n33_n297# a_n269_n200# a_207_n200# a_159_n297#
+ a_63_231# VSUBS
X0 a_n177_n200# a_n225_n297# a_n269_n200# w_n407_n419# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.33 as=0.62 ps=4.62 w=2 l=0.15
X1 a_207_n200# a_159_n297# a_111_n200# w_n407_n419# sky130_fd_pr__pfet_01v8 ad=0.62 pd=4.62 as=0.33 ps=2.33 w=2 l=0.15
X2 a_111_n200# a_63_231# a_15_n200# w_n407_n419# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X3 a_n81_n200# a_n129_231# a_n177_n200# w_n407_n419# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
X4 a_15_n200# a_n33_n297# a_n81_n200# w_n407_n419# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.33 as=0.33 ps=2.33 w=2 l=0.15
C0 a_n33_n297# a_15_n200# 0.01649f
C1 a_111_n200# w_n407_n419# 0.020004f
C2 a_n33_n297# a_n225_n297# 0.025732f
C3 a_n269_n200# a_n177_n200# 0.296004f
C4 a_111_n200# a_159_n297# 0.01649f
C5 a_n81_n200# w_n407_n419# 0.020004f
C6 a_n81_n200# a_n129_231# 0.01649f
C7 a_63_231# a_15_n200# 0.01649f
C8 a_n269_n200# a_n225_n297# 0.01649f
C9 a_111_n200# a_207_n200# 0.296004f
C10 w_n407_n419# a_n129_231# 0.123228f
C11 a_n225_n297# a_n177_n200# 0.01649f
C12 a_n33_n297# a_n81_n200# 0.01649f
C13 a_63_231# a_111_n200# 0.01649f
C14 w_n407_n419# a_159_n297# 0.127948f
C15 a_n33_n297# w_n407_n419# 0.112503f
C16 a_n33_n297# a_n129_231# 0.012606f
C17 a_15_n200# a_111_n200# 0.296004f
C18 w_n407_n419# a_207_n200# 0.14551f
C19 a_n81_n200# a_n177_n200# 0.296004f
C20 a_n33_n297# a_159_n297# 0.025732f
C21 a_n269_n200# w_n407_n419# 0.14551f
C22 a_15_n200# a_n81_n200# 0.296004f
C23 w_n407_n419# a_n177_n200# 0.020004f
C24 a_n129_231# a_n177_n200# 0.01649f
C25 a_63_231# w_n407_n419# 0.123228f
C26 a_159_n297# a_207_n200# 0.01649f
C27 a_63_231# a_n129_231# 0.025732f
C28 a_15_n200# w_n407_n419# 0.020004f
C29 a_n225_n297# w_n407_n419# 0.127948f
C30 a_n225_n297# a_n129_231# 0.012606f
C31 a_63_231# a_159_n297# 0.012606f
C32 a_63_231# a_n33_n297# 0.012606f
C33 a_207_n200# VSUBS 0.092849f
C34 a_111_n200# VSUBS 0.027344f
C35 a_15_n200# VSUBS 0.027344f
C36 a_n81_n200# VSUBS 0.027344f
C37 a_n177_n200# VSUBS 0.027344f
C38 a_n269_n200# VSUBS 0.092849f
C39 a_159_n297# VSUBS 0.061983f
C40 a_n33_n297# VSUBS 0.045346f
C41 a_n225_n297# VSUBS 0.061983f
C42 a_63_231# VSUBS 0.055009f
C43 a_n129_231# VSUBS 0.055009f
C44 w_n407_n419# VSUBS 2.8079f
.ends

.subckt sky130_fd_pr__nfet_01v8_MSLS59 a_n33_n300# a_15_n388# a_n81_322# a_n177_n388#
+ a_159_n300# a_n323_n474# a_n221_n300# a_n129_n300# a_63_n300# a_111_322#
X0 a_159_n300# a_111_322# a_63_n300# a_n323_n474# sky130_fd_pr__nfet_01v8 ad=0.93 pd=6.62 as=0.495 ps=3.33 w=3 l=0.15
X1 a_63_n300# a_15_n388# a_n33_n300# a_n323_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
X2 a_n129_n300# a_n177_n388# a_n221_n300# a_n323_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.93 ps=6.62 w=3 l=0.15
X3 a_n33_n300# a_n81_322# a_n129_n300# a_n323_n474# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=0.15
C0 a_63_n300# a_n33_n300# 0.442473f
C1 a_n177_n388# a_n221_n300# 0.021503f
C2 a_n81_322# a_n33_n300# 0.021503f
C3 a_n177_n388# a_15_n388# 0.02473f
C4 a_n129_n300# a_n81_322# 0.021503f
C5 a_n129_n300# a_n33_n300# 0.442473f
C6 a_159_n300# a_111_322# 0.021503f
C7 a_111_322# a_15_n388# 0.013333f
C8 a_63_n300# a_159_n300# 0.442473f
C9 a_63_n300# a_15_n388# 0.021503f
C10 a_n81_322# a_15_n388# 0.013333f
C11 a_15_n388# a_n33_n300# 0.021503f
C12 a_n129_n300# a_n221_n300# 0.442473f
C13 a_n177_n388# a_n81_322# 0.013333f
C14 a_63_n300# a_111_322# 0.021503f
C15 a_n129_n300# a_n177_n388# 0.021503f
C16 a_n81_322# a_111_322# 0.02473f
C17 a_159_n300# a_n323_n474# 0.340732f
C18 a_63_n300# a_n323_n474# 0.056162f
C19 a_n33_n300# a_n323_n474# 0.056162f
C20 a_n129_n300# a_n323_n474# 0.056162f
C21 a_n221_n300# a_n323_n474# 0.340732f
C22 a_15_n388# a_n323_n474# 0.171561f
C23 a_111_322# a_n323_n474# 0.183396f
C24 a_n177_n388# a_n323_n474# 0.183396f
C25 a_n81_322# a_n323_n474# 0.171561f
.ends

.subckt por_pex VDD Va PAD Vb VSS Vout
Xsky130_fd_pr__res_xhigh_po_1p41_VHK7CU_0 li_8098_8866# VSS VDD sky130_fd_pr__res_xhigh_po_1p41_VHK7CU
XXM12 VDD Vb VDD m1_7502_6058# VSS sky130_fd_pr__pfet_01v8_3HMWVM
Xsky130_fd_pr__res_xhigh_po_1p41_VHK7CU_1 PAD VSS VDD sky130_fd_pr__res_xhigh_po_1p41_VHK7CU
XXM13 x5/A m1_7502_6058# x5/A x5/A m1_7502_6058# VDD x5/A m1_7502_6058# m1_7502_6058#
+ m1_7502_6058# m1_7502_6058# x5/A VDD VDD m1_7502_6058# VDD m1_7502_6058# m1_7502_6058#
+ VDD VDD m1_7502_6058# x5/A VSS sky130_fd_pr__pfet_01v8_PDPE9S
XXM14 VSS VSS Vb Va Va Vb Va Vb VSS Va VSS Va sky130_fd_pr__nfet_01v8_SC2JGL
Xsky130_fd_pr__res_xhigh_po_1p41_VHK7CU_2 x2/A VSS PAD sky130_fd_pr__res_xhigh_po_1p41_VHK7CU
Xx2 x2/A VSS VSS VDD VDD x2/Y sky130_fd_sc_hd__inv_1
XXM15 Va Vb VDD VDD VSS sky130_fd_pr__pfet_01v8_XGSNAL
Xsky130_fd_pr__nfet_01v8_6H2JYD_0 Va x2/Y VSS VSS sky130_fd_pr__nfet_01v8_6H2JYD
XXM16 Vb VDD Va VDD VSS sky130_fd_pr__pfet_01v8_KRS3CJ
Xx5 x5/A x6/Y VSS VSS VDD VDD Vout x5/a_123_47# x5/a_40_47# sky130_fd_sc_hd__and2_0
Xx6 Vb VSS VSS VDD VDD x6/Y sky130_fd_sc_hd__inv_1
XXM3 m1_9068_8792# Va Va Va m1_9068_8792# m1_9068_8792# dw_8516_8522# dw_8516_8522#
+ Va dw_8516_8522# sky130_fd_pr__nfet_01v8_BBNS5R
XXM4 m1_5506_9002# li_5442_5626# m1_5506_9002# li_5442_5626# VSS sky130_fd_pr__pfet_01v8_SKB8VM
XXM5 m1_5484_9862# m1_5506_9002# m1_5506_9002# m1_5484_9862# VSS sky130_fd_pr__pfet_01v8_SKB8VM
XXM6 VDD m1_5484_9862# m1_5484_9862# VDD VSS sky130_fd_pr__pfet_01v8_SKB8VM
XXM7 li_5442_5626# Va li_5442_5626# x2/Y x2/Y Va x2/Y x2/Y x2/Y li_5442_5626# Va Va
+ x2/Y x2/Y li_5442_5626# Va x2/Y li_5442_5626# li_5442_5626# x2/Y Va x2/Y VSS sky130_fd_pr__pfet_01v8_VC5S4W
XXM8 VSS VSS x5/A m1_7502_6058# sky130_fd_pr__nfet_01v8_69TQ3K
XXM9 m1_9068_8792# m1_9068_8792# Va m1_9068_8792# li_8098_8866# li_8098_8866# li_8098_8866#
+ Va Va Va VSS sky130_fd_pr__pfet_01v8_UGNVTG
Xsky130_fd_pr__nfet_01v8_U2JGXT_0 dw_8516_8522# VSS dw_8516_8522# VSS sky130_fd_pr__nfet_01v8_U2JGXT
XXM10 VDD VDD m1_9068_8792# Va VDD m1_9068_8792# Va m1_9068_8792# Va VDD m1_9068_8792#
+ m1_9068_8792# VSS sky130_fd_pr__pfet_01v8_XGS3BL
XXM11 m1_7502_6058# Vb Vb Vb m1_7502_6058# VSS m1_7502_6058# VSS VSS Vb sky130_fd_pr__nfet_01v8_MSLS59
C0 Vb x5/a_123_47# 2.67e-20
C1 m1_8550_8796# Va 0.024032f
C2 dw_8516_8522# w_8708_8772# 1.834764f
C3 VDD VSS 4.040763f
C4 VSS x2/A 0.501536f
C5 VSS Vout 0.021026f
C6 dw_8516_8522# m1_8550_8968# 0.027969f
C7 dw_8516_8522# w_8516_10738# 0.082663f
C8 VSS m1_5484_9862# 0.058502f
C9 li_8098_8866# x5/a_40_47# 9.57e-19
C10 li_8098_8866# dw_8516_8522# 0.476944f
C11 m1_7502_6058# Va 0.033806f
C12 dw_8516_8522# li_5442_5626# 6.54e-19
C13 VSS x6/Y 0.15951f
C14 m1_5506_9002# Va 0.104017f
C15 Vb x5/a_40_47# 0.002779f
C16 VDD w_8708_8772# -6.1e-23
C17 dw_8516_8522# Vb 0.007714f
C18 VDD PAD 0.292979f
C19 PAD x2/A 0.069679f
C20 li_8098_8866# m2_9036_8556# 0.014202f
C21 li_8098_8866# x5/A 9.33e-19
C22 VDD m1_8550_8968# 7.38e-20
C23 Va m2_9036_8622# 0.025635f
C24 m1_7960_6714# Vb 0.046885f
C25 VDD w_8516_10738# 0.005758f
C26 PAD m1_5484_9862# 0.035634f
C27 Vb x5/A 0.040841f
C28 li_8098_8866# VDD 1.148516f
C29 dw_8516_8522# m1_9068_8792# 1.205927f
C30 VSS Va 3.635144f
C31 VDD li_5442_5626# 0.155899f
C32 li_5442_5626# x2/A 0.08617f
C33 li_8098_8866# Vout 0.002292f
C34 VDD Vb 1.56675f
C35 Vb Vout 0.044771f
C36 li_8098_8866# m1_5484_9862# 0.042915f
C37 li_5442_5626# m1_5484_9862# 0.020972f
C38 m1_7502_6058# VSS 1.889269f
C39 m1_7960_6714# x2/Y 0.003322f
C40 li_8098_8866# x6/Y 0.001711f
C41 m1_5506_9002# VSS 0.153436f
C42 x5/a_123_47# x5/A 5.05e-19
C43 VDD m1_9068_8792# 0.889086f
C44 Va w_8708_8772# 0.021672f
C45 Vb x6/Y 0.044227f
C46 Va PAD 0.026236f
C47 m1_8550_8796# m1_8550_8968# 0.014667f
C48 VDD x2/Y 0.137378f
C49 x2/Y x2/A 0.07108f
C50 VDD x5/a_123_47# -2.54e-19
C51 Va m1_8550_8968# 0.002015f
C52 li_8098_8866# m1_8550_8796# 5.99e-19
C53 m1_9068_8792# m1_5484_9862# 0.065313f
C54 Va w_8516_10738# 0.007591f
C55 li_8098_8866# Va 1.384159f
C56 Va li_5442_5626# 2.947124f
C57 m1_7960_6714# dw_8516_8522# 9.09e-21
C58 m1_5506_9002# PAD 0.079987f
C59 dw_8516_8522# m2_9036_8556# 0.008611f
C60 Vb Va 1.474572f
C61 x5/A x5/a_40_47# 0.015036f
C62 x5/a_123_47# x6/Y 0.001168f
C63 VDD x5/a_40_47# 0.012417f
C64 VDD dw_8516_8522# 0.278543f
C65 m1_8550_8796# m1_9068_8792# 0.005121f
C66 li_8098_8866# m1_5506_9002# 0.006542f
C67 x5/a_40_47# Vout 0.001748f
C68 m1_7502_6058# Vb 0.761893f
C69 m1_5506_9002# li_5442_5626# 0.446639f
C70 VSS PAD 0.438805f
C71 Va m1_9068_8792# 1.618831f
C72 VDD m1_7960_6714# 0.087392f
C73 li_8098_8866# m2_9036_8622# 0.010847f
C74 Va x2/Y 1.477496f
C75 VDD m2_9036_8556# 0.001172f
C76 VDD x5/A 2.325278f
C77 x5/a_40_47# x6/Y 0.039015f
C78 x5/A Vout 0.00692f
C79 li_8098_8866# VSS 0.220987f
C80 VSS li_5442_5626# 0.442061f
C81 VDD x2/A 0.344681f
C82 m1_5506_9002# m1_9068_8792# 0.005198f
C83 Vb VSS 1.739453f
C84 VDD Vout 0.082272f
C85 m1_5506_9002# x2/Y 0.050727f
C86 x5/A x6/Y 0.169689f
C87 m1_9068_8792# m2_9036_8622# 0.003458f
C88 dw_8516_8522# m1_8550_8796# 0.01766f
C89 VDD m1_5484_9862# 0.937134f
C90 dw_8516_8522# Va 1.681919f
C91 VDD x6/Y 0.269024f
C92 VSS m1_9068_8792# 0.009944f
C93 Vout x6/Y 0.003725f
C94 PAD li_5442_5626# 0.174135f
C95 VSS x2/Y 1.076192f
C96 m1_7960_6714# Va 0.10714f
C97 x5/a_123_47# VSS 0.001586f
C98 li_8098_8866# m1_8550_8968# 4.97e-19
C99 m2_9036_8556# Va 0.011079f
C100 m1_7502_6058# x5/a_40_47# 0.004315f
C101 x5/A Va 1.24e-19
C102 VDD m1_8550_8796# 7.38e-20
C103 m1_5506_9002# dw_8516_8522# 2.66e-19
C104 m1_7502_6058# m1_7960_6714# 0.011242f
C105 VDD Va 1.908683f
C106 Va x2/A 7.48e-19
C107 m1_9068_8792# w_8708_8772# 0.001356f
C108 li_8098_8866# Vb 0.270498f
C109 m1_7502_6058# x5/A 1.929988f
C110 Vb li_5442_5626# 0.002181f
C111 dw_8516_8522# m2_9036_8622# 0.018145f
C112 x2/Y PAD 3.82e-19
C113 m1_9068_8792# m1_8550_8968# 0.005297f
C114 Va m1_5484_9862# 0.002148f
C115 VSS x5/a_40_47# 0.039655f
C116 VDD m1_7502_6058# 2.158934f
C117 dw_8516_8522# VSS 0.42024f
C118 m1_9068_8792# w_8516_10738# 0.002346f
C119 m2_9036_8556# m2_9036_8622# 0.040517f
C120 Va x6/Y 2.44e-20
C121 m1_7502_6058# Vout 0.031721f
C122 li_8098_8866# m1_9068_8792# 0.637048f
C123 m1_5506_9002# VDD 0.161042f
C124 m1_7960_6714# VSS 0.006795f
C125 Vb m1_9068_8792# 0.033997f
C126 x2/Y li_5442_5626# 1.176716f
C127 VSS x5/A 0.426603f
C128 m1_7502_6058# x6/Y 0.028198f
C129 m1_5506_9002# m1_5484_9862# 0.554574f
C130 Vb x2/Y 0.087483f
C131 m2_9036_8556# 0 0.009013f $ **FLOATING
C132 m2_9036_8622# 0 9.25e-19 $ **FLOATING
C133 m1_7960_6714# 0 0.092041f $ **FLOATING
C134 m1_8550_8796# 0 2.87e-19 $ **FLOATING
C135 m1_8550_8968# 0 0.002438f $ **FLOATING
C136 VSS 0 11.189935f
C137 dw_8516_8522# 0 7.152397f
C138 m1_9068_8792# 0 2.734346f
C139 li_8098_8866# 0 8.171266f
C140 x5/A 0 2.507575f
C141 Va 0 6.359907f
C142 x2/Y 0 2.407521f
C143 li_5442_5626# 0 11.403434f
C144 m1_5484_9862# 0 6.072351f
C145 m1_5506_9002# 0 5.921825f
C146 x6/Y 0 0.293297f
C147 Vout 0 0.285337f
C148 x5/a_40_47# 0 0.230074f
C149 VDD 0 56.14505f
C150 x2/A 0 2.341672f
C151 PAD 0 3.037107f
C152 m1_7502_6058# 0 5.499955f
C153 Vb 0 9.135328f
.ends

