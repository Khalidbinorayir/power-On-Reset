magic
tech sky130A
magscale 1 2
timestamp 1721889469
<< error_p >>
rect -29 8081 29 8087
rect -29 8047 -17 8081
rect -29 8041 29 8047
rect -29 -8047 29 -8041
rect -29 -8081 -17 -8047
rect -29 -8087 29 -8081
<< nwell >>
rect -211 -8219 211 8219
<< pmos >>
rect -15 -8000 15 8000
<< pdiff >>
rect -73 7988 -15 8000
rect -73 -7988 -61 7988
rect -27 -7988 -15 7988
rect -73 -8000 -15 -7988
rect 15 7988 73 8000
rect 15 -7988 27 7988
rect 61 -7988 73 7988
rect 15 -8000 73 -7988
<< pdiffc >>
rect -61 -7988 -27 7988
rect 27 -7988 61 7988
<< nsubdiff >>
rect -175 8149 -79 8183
rect 79 8149 175 8183
rect -175 8087 -141 8149
rect 141 8087 175 8149
rect -175 -8149 -141 -8087
rect 141 -8149 175 -8087
rect -175 -8183 -79 -8149
rect 79 -8183 175 -8149
<< nsubdiffcont >>
rect -79 8149 79 8183
rect -175 -8087 -141 8087
rect 141 -8087 175 8087
rect -79 -8183 79 -8149
<< poly >>
rect -33 8081 33 8097
rect -33 8047 -17 8081
rect 17 8047 33 8081
rect -33 8031 33 8047
rect -15 8000 15 8031
rect -15 -8031 15 -8000
rect -33 -8047 33 -8031
rect -33 -8081 -17 -8047
rect 17 -8081 33 -8047
rect -33 -8097 33 -8081
<< polycont >>
rect -17 8047 17 8081
rect -17 -8081 17 -8047
<< locali >>
rect -175 8149 -79 8183
rect 79 8149 175 8183
rect -175 8087 -141 8149
rect 141 8087 175 8149
rect -33 8047 -17 8081
rect 17 8047 33 8081
rect -61 7988 -27 8004
rect -61 -8004 -27 -7988
rect 27 7988 61 8004
rect 27 -8004 61 -7988
rect -33 -8081 -17 -8047
rect 17 -8081 33 -8047
rect -175 -8149 -141 -8087
rect 141 -8149 175 -8087
rect -175 -8183 -79 -8149
rect 79 -8183 175 -8149
<< viali >>
rect -17 8047 17 8081
rect -61 -7988 -27 7988
rect 27 -7988 61 7988
rect -17 -8081 17 -8047
<< metal1 >>
rect -29 8081 29 8087
rect -29 8047 -17 8081
rect 17 8047 29 8081
rect -29 8041 29 8047
rect -67 7988 -21 8000
rect -67 -7988 -61 7988
rect -27 -7988 -21 7988
rect -67 -8000 -21 -7988
rect 21 7988 67 8000
rect 21 -7988 27 7988
rect 61 -7988 67 7988
rect 21 -8000 67 -7988
rect -29 -8047 29 -8041
rect -29 -8081 -17 -8047
rect 17 -8081 29 -8047
rect -29 -8087 29 -8081
<< properties >>
string FIXED_BBOX -158 -8166 158 8166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 80.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
