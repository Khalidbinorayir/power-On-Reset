magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_p >>
rect -365 881 -307 887
rect -173 881 -115 887
rect 19 881 77 887
rect 211 881 269 887
rect 403 881 461 887
rect -365 847 -353 881
rect -173 847 -161 881
rect 19 847 31 881
rect 211 847 223 881
rect 403 847 415 881
rect -365 841 -307 847
rect -173 841 -115 847
rect 19 841 77 847
rect 211 841 269 847
rect 403 841 461 847
rect -461 -847 -403 -841
rect -269 -847 -211 -841
rect -77 -847 -19 -841
rect 115 -847 173 -841
rect 307 -847 365 -841
rect -461 -881 -449 -847
rect -269 -881 -257 -847
rect -77 -881 -65 -847
rect 115 -881 127 -847
rect 307 -881 319 -847
rect -461 -887 -403 -881
rect -269 -887 -211 -881
rect -77 -887 -19 -881
rect 115 -887 173 -881
rect 307 -887 365 -881
<< nwell >>
rect -647 -1019 647 1019
<< pmos >>
rect -447 -800 -417 800
rect -351 -800 -321 800
rect -255 -800 -225 800
rect -159 -800 -129 800
rect -63 -800 -33 800
rect 33 -800 63 800
rect 129 -800 159 800
rect 225 -800 255 800
rect 321 -800 351 800
rect 417 -800 447 800
<< pdiff >>
rect -509 788 -447 800
rect -509 -788 -497 788
rect -463 -788 -447 788
rect -509 -800 -447 -788
rect -417 788 -351 800
rect -417 -788 -401 788
rect -367 -788 -351 788
rect -417 -800 -351 -788
rect -321 788 -255 800
rect -321 -788 -305 788
rect -271 -788 -255 788
rect -321 -800 -255 -788
rect -225 788 -159 800
rect -225 -788 -209 788
rect -175 -788 -159 788
rect -225 -800 -159 -788
rect -129 788 -63 800
rect -129 -788 -113 788
rect -79 -788 -63 788
rect -129 -800 -63 -788
rect -33 788 33 800
rect -33 -788 -17 788
rect 17 -788 33 788
rect -33 -800 33 -788
rect 63 788 129 800
rect 63 -788 79 788
rect 113 -788 129 788
rect 63 -800 129 -788
rect 159 788 225 800
rect 159 -788 175 788
rect 209 -788 225 788
rect 159 -800 225 -788
rect 255 788 321 800
rect 255 -788 271 788
rect 305 -788 321 788
rect 255 -800 321 -788
rect 351 788 417 800
rect 351 -788 367 788
rect 401 -788 417 788
rect 351 -800 417 -788
rect 447 788 509 800
rect 447 -788 463 788
rect 497 -788 509 788
rect 447 -800 509 -788
<< pdiffc >>
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
<< nsubdiff >>
rect -611 949 -515 983
rect 515 949 611 983
rect -611 887 -577 949
rect 577 887 611 949
rect -611 -949 -577 -887
rect 577 -949 611 -887
rect -611 -983 -515 -949
rect 515 -983 611 -949
<< nsubdiffcont >>
rect -515 949 515 983
rect -611 -887 -577 887
rect 577 -887 611 887
rect -515 -983 515 -949
<< poly >>
rect -369 881 -303 897
rect -369 847 -353 881
rect -319 847 -303 881
rect -369 831 -303 847
rect -177 881 -111 897
rect -177 847 -161 881
rect -127 847 -111 881
rect -177 831 -111 847
rect 15 881 81 897
rect 15 847 31 881
rect 65 847 81 881
rect 15 831 81 847
rect 207 881 273 897
rect 207 847 223 881
rect 257 847 273 881
rect 207 831 273 847
rect 399 881 465 897
rect 399 847 415 881
rect 449 847 465 881
rect 399 831 465 847
rect -447 800 -417 826
rect -351 800 -321 831
rect -255 800 -225 826
rect -159 800 -129 831
rect -63 800 -33 826
rect 33 800 63 831
rect 129 800 159 826
rect 225 800 255 831
rect 321 800 351 826
rect 417 800 447 831
rect -447 -831 -417 -800
rect -351 -826 -321 -800
rect -255 -831 -225 -800
rect -159 -826 -129 -800
rect -63 -831 -33 -800
rect 33 -826 63 -800
rect 129 -831 159 -800
rect 225 -826 255 -800
rect 321 -831 351 -800
rect 417 -826 447 -800
rect -465 -847 -399 -831
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -465 -897 -399 -881
rect -273 -847 -207 -831
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -273 -897 -207 -881
rect -81 -847 -15 -831
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect -81 -897 -15 -881
rect 111 -847 177 -831
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 111 -897 177 -881
rect 303 -847 369 -831
rect 303 -881 319 -847
rect 353 -881 369 -847
rect 303 -897 369 -881
<< polycont >>
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
<< locali >>
rect -611 949 -515 983
rect 515 949 611 983
rect -611 887 -577 949
rect 577 887 611 949
rect -369 847 -353 881
rect -319 847 -303 881
rect -177 847 -161 881
rect -127 847 -111 881
rect 15 847 31 881
rect 65 847 81 881
rect 207 847 223 881
rect 257 847 273 881
rect 399 847 415 881
rect 449 847 465 881
rect -497 788 -463 804
rect -497 -804 -463 -788
rect -401 788 -367 804
rect -401 -804 -367 -788
rect -305 788 -271 804
rect -305 -804 -271 -788
rect -209 788 -175 804
rect -209 -804 -175 -788
rect -113 788 -79 804
rect -113 -804 -79 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 79 788 113 804
rect 79 -804 113 -788
rect 175 788 209 804
rect 175 -804 209 -788
rect 271 788 305 804
rect 271 -804 305 -788
rect 367 788 401 804
rect 367 -804 401 -788
rect 463 788 497 804
rect 463 -804 497 -788
rect -465 -881 -449 -847
rect -415 -881 -399 -847
rect -273 -881 -257 -847
rect -223 -881 -207 -847
rect -81 -881 -65 -847
rect -31 -881 -15 -847
rect 111 -881 127 -847
rect 161 -881 177 -847
rect 303 -881 319 -847
rect 353 -881 369 -847
rect -611 -949 -577 -887
rect 577 -949 611 -887
rect -611 -983 -515 -949
rect 515 -983 611 -949
<< viali >>
rect -353 847 -319 881
rect -161 847 -127 881
rect 31 847 65 881
rect 223 847 257 881
rect 415 847 449 881
rect -497 -788 -463 788
rect -401 -788 -367 788
rect -305 -788 -271 788
rect -209 -788 -175 788
rect -113 -788 -79 788
rect -17 -788 17 788
rect 79 -788 113 788
rect 175 -788 209 788
rect 271 -788 305 788
rect 367 -788 401 788
rect 463 -788 497 788
rect -449 -881 -415 -847
rect -257 -881 -223 -847
rect -65 -881 -31 -847
rect 127 -881 161 -847
rect 319 -881 353 -847
<< metal1 >>
rect -365 881 -307 887
rect -365 847 -353 881
rect -319 847 -307 881
rect -365 841 -307 847
rect -173 881 -115 887
rect -173 847 -161 881
rect -127 847 -115 881
rect -173 841 -115 847
rect 19 881 77 887
rect 19 847 31 881
rect 65 847 77 881
rect 19 841 77 847
rect 211 881 269 887
rect 211 847 223 881
rect 257 847 269 881
rect 211 841 269 847
rect 403 881 461 887
rect 403 847 415 881
rect 449 847 461 881
rect 403 841 461 847
rect -503 788 -457 800
rect -503 -788 -497 788
rect -463 -788 -457 788
rect -503 -800 -457 -788
rect -407 788 -361 800
rect -407 -788 -401 788
rect -367 -788 -361 788
rect -407 -800 -361 -788
rect -311 788 -265 800
rect -311 -788 -305 788
rect -271 -788 -265 788
rect -311 -800 -265 -788
rect -215 788 -169 800
rect -215 -788 -209 788
rect -175 -788 -169 788
rect -215 -800 -169 -788
rect -119 788 -73 800
rect -119 -788 -113 788
rect -79 -788 -73 788
rect -119 -800 -73 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 73 788 119 800
rect 73 -788 79 788
rect 113 -788 119 788
rect 73 -800 119 -788
rect 169 788 215 800
rect 169 -788 175 788
rect 209 -788 215 788
rect 169 -800 215 -788
rect 265 788 311 800
rect 265 -788 271 788
rect 305 -788 311 788
rect 265 -800 311 -788
rect 361 788 407 800
rect 361 -788 367 788
rect 401 -788 407 788
rect 361 -800 407 -788
rect 457 788 503 800
rect 457 -788 463 788
rect 497 -788 503 788
rect 457 -800 503 -788
rect -461 -847 -403 -841
rect -461 -881 -449 -847
rect -415 -881 -403 -847
rect -461 -887 -403 -881
rect -269 -847 -211 -841
rect -269 -881 -257 -847
rect -223 -881 -211 -847
rect -269 -887 -211 -881
rect -77 -847 -19 -841
rect -77 -881 -65 -847
rect -31 -881 -19 -847
rect -77 -887 -19 -881
rect 115 -847 173 -841
rect 115 -881 127 -847
rect 161 -881 173 -847
rect 115 -887 173 -881
rect 307 -847 365 -841
rect 307 -881 319 -847
rect 353 -881 365 -847
rect 307 -887 365 -881
<< properties >>
string FIXED_BBOX -594 -966 594 966
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 0.15 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
