magic
tech sky130A
magscale 1 2
timestamp 1723031900
<< error_p >>
rect -77 972 -19 978
rect 115 972 173 978
rect -77 938 -65 972
rect 115 938 127 972
rect -77 932 -19 938
rect 115 932 173 938
rect -173 -938 -115 -932
rect 19 -938 77 -932
rect -173 -972 -161 -938
rect 19 -972 31 -938
rect -173 -978 -115 -972
rect 19 -978 77 -972
<< pwell >>
rect -359 -1110 359 1110
<< nmos >>
rect -159 -900 -129 900
rect -63 -900 -33 900
rect 33 -900 63 900
rect 129 -900 159 900
<< ndiff >>
rect -221 888 -159 900
rect -221 -888 -209 888
rect -175 -888 -159 888
rect -221 -900 -159 -888
rect -129 888 -63 900
rect -129 -888 -113 888
rect -79 -888 -63 888
rect -129 -900 -63 -888
rect -33 888 33 900
rect -33 -888 -17 888
rect 17 -888 33 888
rect -33 -900 33 -888
rect 63 888 129 900
rect 63 -888 79 888
rect 113 -888 129 888
rect 63 -900 129 -888
rect 159 888 221 900
rect 159 -888 175 888
rect 209 -888 221 888
rect 159 -900 221 -888
<< ndiffc >>
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
<< psubdiff >>
rect -323 1040 -227 1074
rect 227 1040 323 1074
rect -323 978 -289 1040
rect 289 978 323 1040
rect -323 -1040 -289 -978
rect 289 -1040 323 -978
rect -323 -1074 -227 -1040
rect 227 -1074 323 -1040
<< psubdiffcont >>
rect -227 1040 227 1074
rect -323 -978 -289 978
rect 289 -978 323 978
rect -227 -1074 227 -1040
<< poly >>
rect -81 972 -15 988
rect -81 938 -65 972
rect -31 938 -15 972
rect -159 900 -129 926
rect -81 922 -15 938
rect 111 972 177 988
rect 111 938 127 972
rect 161 938 177 972
rect -63 900 -33 922
rect 33 900 63 926
rect 111 922 177 938
rect 129 900 159 922
rect -159 -922 -129 -900
rect -177 -938 -111 -922
rect -63 -926 -33 -900
rect 33 -922 63 -900
rect -177 -972 -161 -938
rect -127 -972 -111 -938
rect -177 -988 -111 -972
rect 15 -938 81 -922
rect 129 -926 159 -900
rect 15 -972 31 -938
rect 65 -972 81 -938
rect 15 -988 81 -972
<< polycont >>
rect -65 938 -31 972
rect 127 938 161 972
rect -161 -972 -127 -938
rect 31 -972 65 -938
<< locali >>
rect -323 1040 -227 1074
rect 227 1040 323 1074
rect -323 978 -289 1040
rect 289 978 323 1040
rect -81 938 -65 972
rect -31 938 -15 972
rect 111 938 127 972
rect 161 938 177 972
rect -209 888 -175 904
rect -209 -904 -175 -888
rect -113 888 -79 904
rect -113 -904 -79 -888
rect -17 888 17 904
rect -17 -904 17 -888
rect 79 888 113 904
rect 79 -904 113 -888
rect 175 888 209 904
rect 175 -904 209 -888
rect -177 -972 -161 -938
rect -127 -972 -111 -938
rect 15 -972 31 -938
rect 65 -972 81 -938
rect -323 -1040 -289 -978
rect 289 -1040 323 -978
rect -323 -1074 -227 -1040
rect 227 -1074 323 -1040
<< viali >>
rect -65 938 -31 972
rect 127 938 161 972
rect -209 -888 -175 888
rect -113 -888 -79 888
rect -17 -888 17 888
rect 79 -888 113 888
rect 175 -888 209 888
rect -161 -972 -127 -938
rect 31 -972 65 -938
<< metal1 >>
rect -77 972 -19 978
rect -77 938 -65 972
rect -31 938 -19 972
rect -77 932 -19 938
rect 115 972 173 978
rect 115 938 127 972
rect 161 938 173 972
rect 115 932 173 938
rect -215 888 -169 900
rect -215 -888 -209 888
rect -175 -888 -169 888
rect -215 -900 -169 -888
rect -119 888 -73 900
rect -119 -888 -113 888
rect -79 -888 -73 888
rect -119 -900 -73 -888
rect -23 888 23 900
rect -23 -888 -17 888
rect 17 -888 23 888
rect -23 -900 23 -888
rect 73 888 119 900
rect 73 -888 79 888
rect 113 -888 119 888
rect 73 -900 119 -888
rect 169 888 215 900
rect 169 -888 175 888
rect 209 -888 215 888
rect 169 -900 215 -888
rect -173 -938 -115 -932
rect -173 -972 -161 -938
rect -127 -972 -115 -938
rect -173 -978 -115 -972
rect 19 -938 77 -932
rect 19 -972 31 -938
rect 65 -972 77 -938
rect 19 -978 77 -972
<< properties >>
string FIXED_BBOX -306 -1057 306 1057
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 9.0 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
