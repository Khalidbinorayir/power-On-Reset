magic
tech sky130A
magscale 1 2
timestamp 1721895348
<< error_p >>
rect 19 672 77 678
rect 19 638 31 672
rect 19 632 77 638
rect -77 -638 -19 -632
rect -77 -672 -65 -638
rect -77 -678 -19 -672
<< pwell >>
rect -263 -810 263 810
<< nmos >>
rect -63 -600 -33 600
rect 33 -600 63 600
<< ndiff >>
rect -125 588 -63 600
rect -125 -588 -113 588
rect -79 -588 -63 588
rect -125 -600 -63 -588
rect -33 588 33 600
rect -33 -588 -17 588
rect 17 -588 33 588
rect -33 -600 33 -588
rect 63 588 125 600
rect 63 -588 79 588
rect 113 -588 125 588
rect 63 -600 125 -588
<< ndiffc >>
rect -113 -588 -79 588
rect -17 -588 17 588
rect 79 -588 113 588
<< psubdiff >>
rect -227 740 -131 774
rect 131 740 227 774
rect -227 678 -193 740
rect 193 678 227 740
rect -227 -740 -193 -678
rect 193 -740 227 -678
rect -227 -774 -131 -740
rect 131 -774 227 -740
<< psubdiffcont >>
rect -131 740 131 774
rect -227 -678 -193 678
rect 193 -678 227 678
rect -131 -774 131 -740
<< poly >>
rect 15 672 81 688
rect 15 638 31 672
rect 65 638 81 672
rect -63 600 -33 626
rect 15 622 81 638
rect 33 600 63 622
rect -63 -622 -33 -600
rect -81 -638 -15 -622
rect 33 -626 63 -600
rect -81 -672 -65 -638
rect -31 -672 -15 -638
rect -81 -688 -15 -672
<< polycont >>
rect 31 638 65 672
rect -65 -672 -31 -638
<< locali >>
rect -227 740 -131 774
rect 131 740 227 774
rect -227 678 -193 740
rect 193 678 227 740
rect 15 638 31 672
rect 65 638 81 672
rect -113 588 -79 604
rect -113 -604 -79 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 79 588 113 604
rect 79 -604 113 -588
rect -81 -672 -65 -638
rect -31 -672 -15 -638
rect -227 -740 -193 -678
rect 193 -740 227 -678
rect -227 -774 -131 -740
rect 131 -774 227 -740
<< viali >>
rect 31 638 65 672
rect -113 -588 -79 588
rect -17 -588 17 588
rect 79 -588 113 588
rect -65 -672 -31 -638
<< metal1 >>
rect 19 672 77 678
rect 19 638 31 672
rect 65 638 77 672
rect 19 632 77 638
rect -119 588 -73 600
rect -119 -588 -113 588
rect -79 -588 -73 588
rect -119 -600 -73 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 73 588 119 600
rect 73 -588 79 588
rect 113 -588 119 588
rect 73 -600 119 -588
rect -77 -638 -19 -632
rect -77 -672 -65 -638
rect -31 -672 -19 -638
rect -77 -678 -19 -672
<< properties >>
string FIXED_BBOX -210 -757 210 757
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 6.0 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
