magic
tech sky130A
magscale 1 2
timestamp 1721889469
<< error_p >>
rect -29 1272 29 1278
rect -29 1238 -17 1272
rect -29 1232 29 1238
rect -29 -1238 29 -1232
rect -29 -1272 -17 -1238
rect -29 -1278 29 -1272
<< pwell >>
rect -211 -1410 211 1410
<< nmos >>
rect -15 -1200 15 1200
<< ndiff >>
rect -73 1188 -15 1200
rect -73 -1188 -61 1188
rect -27 -1188 -15 1188
rect -73 -1200 -15 -1188
rect 15 1188 73 1200
rect 15 -1188 27 1188
rect 61 -1188 73 1188
rect 15 -1200 73 -1188
<< ndiffc >>
rect -61 -1188 -27 1188
rect 27 -1188 61 1188
<< psubdiff >>
rect -175 1340 -79 1374
rect 79 1340 175 1374
rect -175 1278 -141 1340
rect 141 1278 175 1340
rect -175 -1340 -141 -1278
rect 141 -1340 175 -1278
rect -175 -1374 -79 -1340
rect 79 -1374 175 -1340
<< psubdiffcont >>
rect -79 1340 79 1374
rect -175 -1278 -141 1278
rect 141 -1278 175 1278
rect -79 -1374 79 -1340
<< poly >>
rect -33 1272 33 1288
rect -33 1238 -17 1272
rect 17 1238 33 1272
rect -33 1222 33 1238
rect -15 1200 15 1222
rect -15 -1222 15 -1200
rect -33 -1238 33 -1222
rect -33 -1272 -17 -1238
rect 17 -1272 33 -1238
rect -33 -1288 33 -1272
<< polycont >>
rect -17 1238 17 1272
rect -17 -1272 17 -1238
<< locali >>
rect -175 1340 -79 1374
rect 79 1340 175 1374
rect -175 1278 -141 1340
rect 141 1278 175 1340
rect -33 1238 -17 1272
rect 17 1238 33 1272
rect -61 1188 -27 1204
rect -61 -1204 -27 -1188
rect 27 1188 61 1204
rect 27 -1204 61 -1188
rect -33 -1272 -17 -1238
rect 17 -1272 33 -1238
rect -175 -1340 -141 -1278
rect 141 -1340 175 -1278
rect -175 -1374 -79 -1340
rect 79 -1374 175 -1340
<< viali >>
rect -17 1238 17 1272
rect -61 -1188 -27 1188
rect 27 -1188 61 1188
rect -17 -1272 17 -1238
<< metal1 >>
rect -29 1272 29 1278
rect -29 1238 -17 1272
rect 17 1238 29 1272
rect -29 1232 29 1238
rect -67 1188 -21 1200
rect -67 -1188 -61 1188
rect -27 -1188 -21 1188
rect -67 -1200 -21 -1188
rect 21 1188 67 1200
rect 21 -1188 27 1188
rect 61 -1188 67 1188
rect 21 -1200 67 -1188
rect -29 -1238 29 -1232
rect -29 -1272 -17 -1238
rect 17 -1272 29 -1238
rect -29 -1278 29 -1272
<< properties >>
string FIXED_BBOX -158 -1357 158 1357
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 12.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
